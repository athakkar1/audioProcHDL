
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;
library WORK;
USE work.arraypkg.ALL;

package sinewave is
  constant wave : mem := (
to_signed(0, 24), to_signed(12867, 24), to_signed(25735, 24), to_signed(38603, 24), to_signed(51471, 24), to_signed(64339, 24), to_signed(77206, 24), to_signed(90074, 24), to_signed(102941, 24), to_signed(115807, 24), to_signed(128674, 24), to_signed(141540, 24), to_signed(154406, 24), to_signed(167272, 24), to_signed(180137, 24), to_signed(193002, 24), to_signed(205866, 24), to_signed(218730, 24), to_signed(231593, 24), to_signed(244456, 24), to_signed(257318, 24), to_signed(270180, 24), to_signed(283041, 24), to_signed(295901, 24), to_signed(308761, 24), to_signed(321620, 24), to_signed(334478, 24), to_signed(347335, 24), to_signed(360192, 24), to_signed(373047, 24), to_signed(385902, 24), to_signed(398756, 24), to_signed(411609, 24), to_signed(424461, 24), to_signed(437312, 24), to_signed(450162, 24), to_signed(463011, 24), to_signed(475859, 24), to_signed(488705, 24), to_signed(501551, 24), to_signed(514395, 24), to_signed(527238, 24), to_signed(540080, 24), to_signed(552921, 24), to_signed(565760, 24), to_signed(578598, 24), to_signed(591435, 24), to_signed(604270, 24), to_signed(617104, 24), to_signed(629936, 24), to_signed(642767, 24), to_signed(655596, 24), to_signed(668424, 24), to_signed(681250, 24), to_signed(694075, 24), to_signed(706898, 24), to_signed(719720, 24), to_signed(732539, 24), to_signed(745357, 24), to_signed(758173, 24), to_signed(770988, 24), to_signed(783800, 24), to_signed(796611, 24), to_signed(809420, 24), to_signed(822227, 24), to_signed(835032, 24), to_signed(847835, 24), to_signed(860636, 24), to_signed(873435, 24), to_signed(886232, 24), to_signed(899027, 24), to_signed(911820, 24), to_signed(924610, 24), to_signed(937399, 24), to_signed(950185, 24), to_signed(962969, 24), to_signed(975751, 24), to_signed(988530, 24), to_signed(1001307, 24), to_signed(1014082, 24), to_signed(1026855, 24), to_signed(1039625, 24), to_signed(1052392, 24), to_signed(1065157, 24), to_signed(1077920, 24), to_signed(1090680, 24), to_signed(1103437, 24), to_signed(1116192, 24), to_signed(1128944, 24), to_signed(1141694, 24), to_signed(1154441, 24), to_signed(1167185, 24), to_signed(1179926, 24), to_signed(1192665, 24), to_signed(1205401, 24), to_signed(1218134, 24), to_signed(1230864, 24), to_signed(1243591, 24), to_signed(1256315, 24), to_signed(1269037, 24), to_signed(1281755, 24), to_signed(1294471, 24), to_signed(1307183, 24), to_signed(1319892, 24), to_signed(1332598, 24), to_signed(1345301, 24), to_signed(1358001, 24), to_signed(1370698, 24), to_signed(1383391, 24), to_signed(1396081, 24), to_signed(1408768, 24), to_signed(1421452, 24), to_signed(1434132, 24), to_signed(1446809, 24), to_signed(1459482, 24), to_signed(1472152, 24), to_signed(1484819, 24), to_signed(1497482, 24), to_signed(1510141, 24), to_signed(1522797, 24), to_signed(1535449, 24), to_signed(1548098, 24), to_signed(1560743, 24), to_signed(1573385, 24), to_signed(1586022, 24), to_signed(1598656, 24), to_signed(1611287, 24), to_signed(1623913, 24), to_signed(1636536, 24), to_signed(1649155, 24), to_signed(1661769, 24), to_signed(1674380, 24), to_signed(1686987, 24), to_signed(1699591, 24), to_signed(1712190, 24), to_signed(1724785, 24), to_signed(1737376, 24), to_signed(1749963, 24), to_signed(1762545, 24), to_signed(1775124, 24), to_signed(1787698, 24), to_signed(1800269, 24), to_signed(1812835, 24), to_signed(1825396, 24), to_signed(1837954, 24), to_signed(1850507, 24), to_signed(1863056, 24), to_signed(1875600, 24), to_signed(1888140, 24), to_signed(1900676, 24), to_signed(1913207, 24), to_signed(1925733, 24), to_signed(1938255, 24), to_signed(1950773, 24), to_signed(1963286, 24), to_signed(1975794, 24), to_signed(1988298, 24), to_signed(2000797, 24), to_signed(2013291, 24), to_signed(2025780, 24), to_signed(2038265, 24), to_signed(2050745, 24), to_signed(2063220, 24), to_signed(2075690, 24), to_signed(2088156, 24), to_signed(2100616, 24), to_signed(2113072, 24), to_signed(2125522, 24), to_signed(2137968, 24), to_signed(2150408, 24), to_signed(2162844, 24), to_signed(2175274, 24), to_signed(2187699, 24), to_signed(2200119, 24), to_signed(2212534, 24), to_signed(2224944, 24), to_signed(2237348, 24), to_signed(2249747, 24), to_signed(2262141, 24), to_signed(2274530, 24), to_signed(2286913, 24), to_signed(2299291, 24), to_signed(2311663, 24), to_signed(2324030, 24), to_signed(2336392, 24), to_signed(2348748, 24), to_signed(2361099, 24), to_signed(2373443, 24), to_signed(2385783, 24), to_signed(2398117, 24), to_signed(2410445, 24), to_signed(2422767, 24), to_signed(2435084, 24), to_signed(2447395, 24), to_signed(2459700, 24), to_signed(2472000, 24), to_signed(2484293, 24), to_signed(2496581, 24), to_signed(2508863, 24), to_signed(2521139, 24), to_signed(2533409, 24), to_signed(2545673, 24), to_signed(2557931, 24), to_signed(2570183, 24), to_signed(2582429, 24), to_signed(2594669, 24), to_signed(2606903, 24), to_signed(2619131, 24), to_signed(2631353, 24), to_signed(2643568, 24), to_signed(2655777, 24), to_signed(2667980, 24), to_signed(2680177, 24), to_signed(2692367, 24), to_signed(2704551, 24), to_signed(2716729, 24), to_signed(2728900, 24), to_signed(2741065, 24), to_signed(2753223, 24), to_signed(2765375, 24), to_signed(2777521, 24), to_signed(2789659, 24), to_signed(2801792, 24), to_signed(2813917, 24), to_signed(2826036, 24), to_signed(2838149, 24), to_signed(2850255, 24), to_signed(2862354, 24), to_signed(2874446, 24), to_signed(2886531, 24), to_signed(2898610, 24), to_signed(2910682, 24), to_signed(2922747, 24), to_signed(2934805, 24), to_signed(2946857, 24), to_signed(2958901, 24), to_signed(2970938, 24), to_signed(2982969, 24), to_signed(2994992, 24), to_signed(3007009, 24), to_signed(3019018, 24), to_signed(3031020, 24), to_signed(3043015, 24), to_signed(3055003, 24), to_signed(3066984, 24), to_signed(3078957, 24), to_signed(3090923, 24), to_signed(3102882, 24), to_signed(3114834, 24), to_signed(3126778, 24), to_signed(3138715, 24), to_signed(3150645, 24), to_signed(3162567, 24), to_signed(3174482, 24), to_signed(3186389, 24), to_signed(3198289, 24), to_signed(3210181, 24), to_signed(3222065, 24), to_signed(3233943, 24), to_signed(3245812, 24), to_signed(3257674, 24), to_signed(3269528, 24), to_signed(3281375, 24), to_signed(3293213, 24), to_signed(3305044, 24), to_signed(3316868, 24), to_signed(3328683, 24), to_signed(3340491, 24), to_signed(3352290, 24), to_signed(3364082, 24), to_signed(3375866, 24), to_signed(3387642, 24), to_signed(3399410, 24), to_signed(3411170, 24), to_signed(3422922, 24), to_signed(3434666, 24), to_signed(3446402, 24), to_signed(3458130, 24), to_signed(3469849, 24), to_signed(3481561, 24), to_signed(3493264, 24), to_signed(3504959, 24), to_signed(3516646, 24), to_signed(3528324, 24), to_signed(3539994, 24), to_signed(3551656, 24), to_signed(3563310, 24), to_signed(3574955, 24), to_signed(3586592, 24), to_signed(3598220, 24), to_signed(3609840, 24), to_signed(3621451, 24), to_signed(3633054, 24), to_signed(3644648, 24), to_signed(3656234, 24), to_signed(3667811, 24), to_signed(3679379, 24), to_signed(3690939, 24), to_signed(3702490, 24), to_signed(3714032, 24), to_signed(3725566, 24), to_signed(3737091, 24), to_signed(3748607, 24), to_signed(3760114, 24), to_signed(3771613, 24), to_signed(3783102, 24), to_signed(3794583, 24), to_signed(3806055, 24), to_signed(3817517, 24), to_signed(3828971, 24), to_signed(3840416, 24), to_signed(3851852, 24), to_signed(3863278, 24), to_signed(3874696, 24), to_signed(3886104, 24), to_signed(3897504, 24), to_signed(3908894, 24), to_signed(3920275, 24), to_signed(3931646, 24), to_signed(3943009, 24), to_signed(3954362, 24), to_signed(3965706, 24), to_signed(3977040, 24), to_signed(3988366, 24), to_signed(3999681, 24), to_signed(4010988, 24), to_signed(4022285, 24), to_signed(4033572, 24), to_signed(4044850, 24), to_signed(4056119, 24), to_signed(4067378, 24), to_signed(4078627, 24), to_signed(4089867, 24), to_signed(4101097, 24), to_signed(4112317, 24), to_signed(4123528, 24), to_signed(4134729, 24), to_signed(4145921, 24), to_signed(4157102, 24), to_signed(4168274, 24), to_signed(4179436, 24), to_signed(4190588, 24), to_signed(4201731, 24), to_signed(4212863, 24), to_signed(4223986, 24), to_signed(4235098, 24), to_signed(4246201, 24), to_signed(4257293, 24), to_signed(4268376, 24), to_signed(4279449, 24), to_signed(4290511, 24), to_signed(4301564, 24), to_signed(4312606, 24), to_signed(4323638, 24), to_signed(4334660, 24), to_signed(4345672, 24), to_signed(4356673, 24), to_signed(4367665, 24), to_signed(4378646, 24), to_signed(4389616, 24), to_signed(4400577, 24), to_signed(4411527, 24), to_signed(4422466, 24), to_signed(4433396, 24), to_signed(4444314, 24), to_signed(4455223, 24), to_signed(4466121, 24), to_signed(4477008, 24), to_signed(4487885, 24), to_signed(4498751, 24), to_signed(4509607, 24), to_signed(4520452, 24), to_signed(4531286, 24), to_signed(4542110, 24), to_signed(4552923, 24), to_signed(4563725, 24), to_signed(4574517, 24), to_signed(4585298, 24), to_signed(4596068, 24), to_signed(4606827, 24), to_signed(4617576, 24), to_signed(4628313, 24), to_signed(4639040, 24), to_signed(4649756, 24), to_signed(4660460, 24), to_signed(4671154, 24), to_signed(4681837, 24), to_signed(4692509, 24), to_signed(4703170, 24), to_signed(4713819, 24), to_signed(4724458, 24), to_signed(4735086, 24), to_signed(4745702, 24), to_signed(4756307, 24), to_signed(4766901, 24), to_signed(4777484, 24), to_signed(4788055, 24), to_signed(4798616, 24), to_signed(4809165, 24), to_signed(4819702, 24), to_signed(4830229, 24), to_signed(4840744, 24), to_signed(4851247, 24), to_signed(4861739, 24), to_signed(4872220, 24), to_signed(4882689, 24), to_signed(4893147, 24), to_signed(4903593, 24), to_signed(4914028, 24), to_signed(4924451, 24), to_signed(4934863, 24), to_signed(4945263, 24), to_signed(4955651, 24), to_signed(4966028, 24), to_signed(4976393, 24), to_signed(4986746, 24), to_signed(4997087, 24), to_signed(5007417, 24), to_signed(5017735, 24), to_signed(5028041, 24), to_signed(5038336, 24), to_signed(5048618, 24), to_signed(5058889, 24), to_signed(5069147, 24), to_signed(5079394, 24), to_signed(5089629, 24), to_signed(5099852, 24), to_signed(5110063, 24), to_signed(5120262, 24), to_signed(5130448, 24), to_signed(5140623, 24), to_signed(5150786, 24), to_signed(5160936, 24), to_signed(5171074, 24), to_signed(5181201, 24), to_signed(5191315, 24), to_signed(5201416, 24), to_signed(5211506, 24), to_signed(5221583, 24), to_signed(5231648, 24), to_signed(5241701, 24), to_signed(5251741, 24), to_signed(5261769, 24), to_signed(5271785, 24), to_signed(5281788, 24), to_signed(5291779, 24), to_signed(5301757, 24), to_signed(5311723, 24), to_signed(5321676, 24), to_signed(5331617, 24), to_signed(5341545, 24), to_signed(5351461, 24), to_signed(5361364, 24), to_signed(5371254, 24), to_signed(5381132, 24), to_signed(5390997, 24), to_signed(5400850, 24), to_signed(5410690, 24), to_signed(5420517, 24), to_signed(5430331, 24), to_signed(5440133, 24), to_signed(5449921, 24), to_signed(5459697, 24), to_signed(5469460, 24), to_signed(5479210, 24), to_signed(5488948, 24), to_signed(5498672, 24), to_signed(5508384, 24), to_signed(5518082, 24), to_signed(5527767, 24), to_signed(5537440, 24), to_signed(5547099, 24), to_signed(5556746, 24), to_signed(5566379, 24), to_signed(5575999, 24), to_signed(5585606, 24), to_signed(5595200, 24), to_signed(5604781, 24), to_signed(5614349, 24), to_signed(5623903, 24), to_signed(5633444, 24), to_signed(5642972, 24), to_signed(5652487, 24), to_signed(5661988, 24), to_signed(5671476, 24), to_signed(5680951, 24), to_signed(5690412, 24), to_signed(5699860, 24), to_signed(5709294, 24), to_signed(5718716, 24), to_signed(5728123, 24), to_signed(5737517, 24), to_signed(5746898, 24), to_signed(5756265, 24), to_signed(5765618, 24), to_signed(5774958, 24), to_signed(5784285, 24), to_signed(5793598, 24), to_signed(5802897, 24), to_signed(5812182, 24), to_signed(5821454, 24), to_signed(5830712, 24), to_signed(5839957, 24), to_signed(5849187, 24), to_signed(5858404, 24), to_signed(5867607, 24), to_signed(5876796, 24), to_signed(5885972, 24), to_signed(5895134, 24), to_signed(5904281, 24), to_signed(5913415, 24), to_signed(5922535, 24), to_signed(5931641, 24), to_signed(5940733, 24), to_signed(5949811, 24), to_signed(5958875, 24), to_signed(5967925, 24), to_signed(5976961, 24), to_signed(5985983, 24), to_signed(5994991, 24), to_signed(6003985, 24), to_signed(6012964, 24), to_signed(6021930, 24), to_signed(6030881, 24), to_signed(6039818, 24), to_signed(6048741, 24), to_signed(6057650, 24), to_signed(6066544, 24), to_signed(6075424, 24), to_signed(6084290, 24), to_signed(6093142, 24), to_signed(6101979, 24), to_signed(6110802, 24), to_signed(6119610, 24), to_signed(6128404, 24), to_signed(6137184, 24), to_signed(6145949, 24), to_signed(6154700, 24), to_signed(6163436, 24), to_signed(6172158, 24), to_signed(6180865, 24), to_signed(6189558, 24), to_signed(6198236, 24), to_signed(6206899, 24), to_signed(6215548, 24), to_signed(6224182, 24), to_signed(6232802, 24), to_signed(6241407, 24), to_signed(6249997, 24), to_signed(6258573, 24), to_signed(6267134, 24), to_signed(6275680, 24), to_signed(6284211, 24), to_signed(6292728, 24), to_signed(6301229, 24), to_signed(6309716, 24), to_signed(6318188, 24), to_signed(6326646, 24), to_signed(6335088, 24), to_signed(6343515, 24), to_signed(6351928, 24), to_signed(6360325, 24), to_signed(6368708, 24), to_signed(6377075, 24), to_signed(6385428, 24), to_signed(6393765, 24), to_signed(6402088, 24), to_signed(6410395, 24), to_signed(6418688, 24), to_signed(6426965, 24), to_signed(6435227, 24), to_signed(6443474, 24), to_signed(6451706, 24), to_signed(6459923, 24), to_signed(6468124, 24), to_signed(6476310, 24), to_signed(6484481, 24), to_signed(6492637, 24), to_signed(6500777, 24), to_signed(6508902, 24), to_signed(6517012, 24), to_signed(6525107, 24), to_signed(6533186, 24), to_signed(6541250, 24), to_signed(6549298, 24), to_signed(6557331, 24), to_signed(6565349, 24), to_signed(6573351, 24), to_signed(6581337, 24), to_signed(6589308, 24), to_signed(6597264, 24), to_signed(6605204, 24), to_signed(6613129, 24), to_signed(6621038, 24), to_signed(6628931, 24), to_signed(6636809, 24), to_signed(6644671, 24), to_signed(6652518, 24), to_signed(6660349, 24), to_signed(6668164, 24), to_signed(6675963, 24), to_signed(6683747, 24), to_signed(6691515, 24), to_signed(6699268, 24), to_signed(6707004, 24), to_signed(6714725, 24), to_signed(6722430, 24), to_signed(6730119, 24), to_signed(6737793, 24), to_signed(6745450, 24), to_signed(6753092, 24), to_signed(6760718, 24), to_signed(6768327, 24), to_signed(6775921, 24), to_signed(6783499, 24), to_signed(6791061, 24), to_signed(6798607, 24), to_signed(6806137, 24), to_signed(6813651, 24), to_signed(6821149, 24), to_signed(6828631, 24), to_signed(6836097, 24), to_signed(6843547, 24), to_signed(6850980, 24), to_signed(6858398, 24), to_signed(6865799, 24), to_signed(6873185, 24), to_signed(6880554, 24), to_signed(6887907, 24), to_signed(6895243, 24), to_signed(6902564, 24), to_signed(6909868, 24), to_signed(6917156, 24), to_signed(6924428, 24), to_signed(6931683, 24), to_signed(6938922, 24), to_signed(6946145, 24), to_signed(6953351, 24), to_signed(6960541, 24), to_signed(6967715, 24), to_signed(6974872, 24), to_signed(6982013, 24), to_signed(6989137, 24), to_signed(6996245, 24), to_signed(7003337, 24), to_signed(7010412, 24), to_signed(7017470, 24), to_signed(7024512, 24), to_signed(7031538, 24), to_signed(7038547, 24), to_signed(7045539, 24), to_signed(7052515, 24), to_signed(7059474, 24), to_signed(7066417, 24), to_signed(7073343, 24), to_signed(7080252, 24), to_signed(7087145, 24), to_signed(7094021, 24), to_signed(7100880, 24), to_signed(7107723, 24), to_signed(7114549, 24), to_signed(7121358, 24), to_signed(7128150, 24), to_signed(7134926, 24), to_signed(7141684, 24), to_signed(7148426, 24), to_signed(7155152, 24), to_signed(7161860, 24), to_signed(7168551, 24), to_signed(7175226, 24), to_signed(7181884, 24), to_signed(7188525, 24), to_signed(7195149, 24), to_signed(7201756, 24), to_signed(7208346, 24), to_signed(7214919, 24), to_signed(7221475, 24), to_signed(7228014, 24), to_signed(7234536, 24), to_signed(7241041, 24), to_signed(7247529, 24), to_signed(7254000, 24), to_signed(7260454, 24), to_signed(7266891, 24), to_signed(7273311, 24), to_signed(7279713, 24), to_signed(7286099, 24), to_signed(7292467, 24), to_signed(7298818, 24), to_signed(7305152, 24), to_signed(7311469, 24), to_signed(7317769, 24), to_signed(7324051, 24), to_signed(7330316, 24), to_signed(7336564, 24), to_signed(7342795, 24), to_signed(7349008, 24), to_signed(7355204, 24), to_signed(7361383, 24), to_signed(7367544, 24), to_signed(7373688, 24), to_signed(7379815, 24), to_signed(7385925, 24), to_signed(7392017, 24), to_signed(7398091, 24), to_signed(7404148, 24), to_signed(7410188, 24), to_signed(7416211, 24), to_signed(7422216, 24), to_signed(7428203, 24), to_signed(7434173, 24), to_signed(7440125, 24), to_signed(7446060, 24), to_signed(7451978, 24), to_signed(7457878, 24), to_signed(7463760, 24), to_signed(7469625, 24), to_signed(7475472, 24), to_signed(7481302, 24), to_signed(7487114, 24), to_signed(7492908, 24), to_signed(7498685, 24), to_signed(7504444, 24), to_signed(7510185, 24), to_signed(7515909, 24), to_signed(7521615, 24), to_signed(7527304, 24), to_signed(7532974, 24), to_signed(7538627, 24), to_signed(7544263, 24), to_signed(7549880, 24), to_signed(7555480, 24), to_signed(7561062, 24), to_signed(7566626, 24), to_signed(7572172, 24), to_signed(7577701, 24), to_signed(7583211, 24), to_signed(7588704, 24), to_signed(7594179, 24), to_signed(7599636, 24), to_signed(7605075, 24), to_signed(7610497, 24), to_signed(7615900, 24), to_signed(7621286, 24), to_signed(7626653, 24), to_signed(7632003, 24), to_signed(7637335, 24), to_signed(7642648, 24), to_signed(7647944, 24), to_signed(7653222, 24), to_signed(7658481, 24), to_signed(7663723, 24), to_signed(7668947, 24), to_signed(7674152, 24), to_signed(7679340, 24), to_signed(7684509, 24), to_signed(7689661, 24), to_signed(7694794, 24), to_signed(7699909, 24), to_signed(7705006, 24), to_signed(7710085, 24), to_signed(7715146, 24), to_signed(7720189, 24), to_signed(7725213, 24), to_signed(7730220, 24), to_signed(7735208, 24), to_signed(7740178, 24), to_signed(7745129, 24), to_signed(7750063, 24), to_signed(7754978, 24), to_signed(7759875, 24), to_signed(7764754, 24), to_signed(7769614, 24), to_signed(7774456, 24), to_signed(7779280, 24), to_signed(7784086, 24), to_signed(7788873, 24), to_signed(7793642, 24), to_signed(7798393, 24), to_signed(7803125, 24), to_signed(7807839, 24), to_signed(7812534, 24), to_signed(7817211, 24), to_signed(7821870, 24), to_signed(7826510, 24), to_signed(7831132, 24), to_signed(7835736, 24), to_signed(7840321, 24), to_signed(7844887, 24), to_signed(7849436, 24), to_signed(7853965, 24), to_signed(7858476, 24), to_signed(7862969, 24), to_signed(7867443, 24), to_signed(7871899, 24), to_signed(7876336, 24), to_signed(7880755, 24), to_signed(7885155, 24), to_signed(7889536, 24), to_signed(7893899, 24), to_signed(7898244, 24), to_signed(7902569, 24), to_signed(7906877, 24), to_signed(7911165, 24), to_signed(7915435, 24), to_signed(7919686, 24), to_signed(7923919, 24), to_signed(7928133, 24), to_signed(7932329, 24), to_signed(7936505, 24), to_signed(7940663, 24), to_signed(7944803, 24), to_signed(7948924, 24), to_signed(7953026, 24), to_signed(7957109, 24), to_signed(7961173, 24), to_signed(7965219, 24), to_signed(7969246, 24), to_signed(7973255, 24), to_signed(7977244, 24), to_signed(7981215, 24), to_signed(7985167, 24), to_signed(7989100, 24), to_signed(7993015, 24), to_signed(7996910, 24), to_signed(8000787, 24), to_signed(8004645, 24), to_signed(8008484, 24), to_signed(8012304, 24), to_signed(8016106, 24), to_signed(8019888, 24), to_signed(8023652, 24), to_signed(8027397, 24), to_signed(8031123, 24), to_signed(8034830, 24), to_signed(8038518, 24), to_signed(8042187, 24), to_signed(8045837, 24), to_signed(8049469, 24), to_signed(8053081, 24), to_signed(8056675, 24), to_signed(8060249, 24), to_signed(8063805, 24), to_signed(8067341, 24), to_signed(8070859, 24), to_signed(8074357, 24), to_signed(8077837, 24), to_signed(8081298, 24), to_signed(8084739, 24), to_signed(8088162, 24), to_signed(8091565, 24), to_signed(8094950, 24), to_signed(8098315, 24), to_signed(8101661, 24), to_signed(8104989, 24), to_signed(8108297, 24), to_signed(8111586, 24), to_signed(8114856, 24), to_signed(8118107, 24), to_signed(8121339, 24), to_signed(8124552, 24), to_signed(8127745, 24), to_signed(8130920, 24), to_signed(8134075, 24), to_signed(8137211, 24), to_signed(8140329, 24), to_signed(8143426, 24), to_signed(8146505, 24), to_signed(8149565, 24), to_signed(8152605, 24), to_signed(8155626, 24), to_signed(8158629, 24), to_signed(8161611, 24), to_signed(8164575, 24), to_signed(8167519, 24), to_signed(8170445, 24), to_signed(8173351, 24), to_signed(8176237, 24), to_signed(8179105, 24), to_signed(8181953, 24), to_signed(8184782, 24), to_signed(8187592, 24), to_signed(8190382, 24), to_signed(8193154, 24), to_signed(8195906, 24), to_signed(8198638, 24), to_signed(8201352, 24), to_signed(8204046, 24), to_signed(8206720, 24), to_signed(8209376, 24), to_signed(8212012, 24), to_signed(8214629, 24), to_signed(8217226, 24), to_signed(8219804, 24), to_signed(8222363, 24), to_signed(8224903, 24), to_signed(8227423, 24), to_signed(8229923, 24), to_signed(8232405, 24), to_signed(8234867, 24), to_signed(8237309, 24), to_signed(8239733, 24), to_signed(8242137, 24), to_signed(8244521, 24), to_signed(8246886, 24), to_signed(8249232, 24), to_signed(8251558, 24), to_signed(8253865, 24), to_signed(8256152, 24), to_signed(8258420, 24), to_signed(8260669, 24), to_signed(8262898, 24), to_signed(8265107, 24), to_signed(8267298, 24), to_signed(8269468, 24), to_signed(8271620, 24), to_signed(8273751, 24), to_signed(8275864, 24), to_signed(8277957, 24), to_signed(8280030, 24), to_signed(8282084, 24), to_signed(8284119, 24), to_signed(8286133, 24), to_signed(8288129, 24), to_signed(8290105, 24), to_signed(8292061, 24), to_signed(8293998, 24), to_signed(8295916, 24), to_signed(8297813, 24), to_signed(8299692, 24), to_signed(8301551, 24), to_signed(8303390, 24), to_signed(8305210, 24), to_signed(8307010, 24), to_signed(8308791, 24), to_signed(8310552, 24), to_signed(8312293, 24), to_signed(8314015, 24), to_signed(8315718, 24), to_signed(8317401, 24), to_signed(8319064, 24), to_signed(8320708, 24), to_signed(8322332, 24), to_signed(8323936, 24), to_signed(8325521, 24), to_signed(8327087, 24), to_signed(8328632, 24), to_signed(8330159, 24), to_signed(8331665, 24), to_signed(8333152, 24), to_signed(8334620, 24), to_signed(8336067, 24), to_signed(8337495, 24), to_signed(8338904, 24), to_signed(8340293, 24), to_signed(8341662, 24), to_signed(8343012, 24), to_signed(8344342, 24), to_signed(8345652, 24), to_signed(8346943, 24), to_signed(8348214, 24), to_signed(8349466, 24), to_signed(8350697, 24), to_signed(8351909, 24), to_signed(8353102, 24), to_signed(8354275, 24), to_signed(8355428, 24), to_signed(8356562, 24), to_signed(8357675, 24), to_signed(8358770, 24), to_signed(8359844, 24), to_signed(8360899, 24), to_signed(8361934, 24), to_signed(8362950, 24), to_signed(8363946, 24), to_signed(8364922, 24), to_signed(8365878, 24), to_signed(8366815, 24), to_signed(8367732, 24), to_signed(8368629, 24), to_signed(8369507, 24), to_signed(8370365, 24), to_signed(8371204, 24), to_signed(8372022, 24), to_signed(8372821, 24), to_signed(8373600, 24), to_signed(8374360, 24), to_signed(8375100, 24), to_signed(8375820, 24), to_signed(8376520, 24), to_signed(8377201, 24), to_signed(8377862, 24), to_signed(8378503, 24), to_signed(8379125, 24), to_signed(8379726, 24), to_signed(8380309, 24), to_signed(8380871, 24), to_signed(8381414, 24), to_signed(8381937, 24), to_signed(8382440, 24), to_signed(8382923, 24), to_signed(8383387, 24), to_signed(8383831, 24), to_signed(8384255, 24), to_signed(8384660, 24), to_signed(8385045, 24), to_signed(8385410, 24), to_signed(8385755, 24), to_signed(8386081, 24), to_signed(8386387, 24), to_signed(8386673, 24), to_signed(8386940, 24), to_signed(8387186, 24), to_signed(8387413, 24), to_signed(8387621, 24), to_signed(8387808, 24), to_signed(8387976, 24), to_signed(8388124, 24), to_signed(8388252, 24), to_signed(8388361, 24), to_signed(8388450, 24), to_signed(8388519, 24), to_signed(8388568, 24), to_signed(8388598, 24), to_signed(8388608, 24), to_signed(8388598, 24), to_signed(8388568, 24), to_signed(8388519, 24), to_signed(8388450, 24), to_signed(8388361, 24), to_signed(8388252, 24), to_signed(8388124, 24), to_signed(8387976, 24), to_signed(8387808, 24), to_signed(8387621, 24), to_signed(8387413, 24), to_signed(8387186, 24), to_signed(8386940, 24), to_signed(8386673, 24), to_signed(8386387, 24), to_signed(8386081, 24), to_signed(8385755, 24), to_signed(8385410, 24), to_signed(8385045, 24), to_signed(8384660, 24), to_signed(8384255, 24), to_signed(8383831, 24), to_signed(8383387, 24), to_signed(8382923, 24), to_signed(8382440, 24), to_signed(8381937, 24), to_signed(8381414, 24), to_signed(8380871, 24), to_signed(8380309, 24), to_signed(8379726, 24), to_signed(8379125, 24), to_signed(8378503, 24), to_signed(8377862, 24), to_signed(8377201, 24), to_signed(8376520, 24), to_signed(8375820, 24), to_signed(8375100, 24), to_signed(8374360, 24), to_signed(8373600, 24), to_signed(8372821, 24), to_signed(8372022, 24), to_signed(8371204, 24), to_signed(8370365, 24), to_signed(8369507, 24), to_signed(8368629, 24), to_signed(8367732, 24), to_signed(8366815, 24), to_signed(8365878, 24), to_signed(8364922, 24), to_signed(8363946, 24), to_signed(8362950, 24), to_signed(8361934, 24), to_signed(8360899, 24), to_signed(8359844, 24), to_signed(8358770, 24), to_signed(8357675, 24), to_signed(8356562, 24), to_signed(8355428, 24), to_signed(8354275, 24), to_signed(8353102, 24), to_signed(8351909, 24), to_signed(8350697, 24), to_signed(8349466, 24), to_signed(8348214, 24), to_signed(8346943, 24), to_signed(8345652, 24), to_signed(8344342, 24), to_signed(8343012, 24), to_signed(8341662, 24), to_signed(8340293, 24), to_signed(8338904, 24), to_signed(8337495, 24), to_signed(8336067, 24), to_signed(8334620, 24), to_signed(8333152, 24), to_signed(8331665, 24), to_signed(8330159, 24), to_signed(8328632, 24), to_signed(8327087, 24), to_signed(8325521, 24), to_signed(8323936, 24), to_signed(8322332, 24), to_signed(8320708, 24), to_signed(8319064, 24), to_signed(8317401, 24), to_signed(8315718, 24), to_signed(8314015, 24), to_signed(8312293, 24), to_signed(8310552, 24), to_signed(8308791, 24), to_signed(8307010, 24), to_signed(8305210, 24), to_signed(8303390, 24), to_signed(8301551, 24), to_signed(8299692, 24), to_signed(8297813, 24), to_signed(8295916, 24), to_signed(8293998, 24), to_signed(8292061, 24), to_signed(8290105, 24), to_signed(8288129, 24), to_signed(8286133, 24), to_signed(8284119, 24), to_signed(8282084, 24), to_signed(8280030, 24), to_signed(8277957, 24), to_signed(8275864, 24), to_signed(8273751, 24), to_signed(8271620, 24), to_signed(8269468, 24), to_signed(8267298, 24), to_signed(8265107, 24), to_signed(8262898, 24), to_signed(8260669, 24), to_signed(8258420, 24), to_signed(8256152, 24), to_signed(8253865, 24), to_signed(8251558, 24), to_signed(8249232, 24), to_signed(8246886, 24), to_signed(8244521, 24), to_signed(8242137, 24), to_signed(8239733, 24), to_signed(8237309, 24), to_signed(8234867, 24), to_signed(8232405, 24), to_signed(8229923, 24), to_signed(8227423, 24), to_signed(8224903, 24), to_signed(8222363, 24), to_signed(8219804, 24), to_signed(8217226, 24), to_signed(8214629, 24), to_signed(8212012, 24), to_signed(8209376, 24), to_signed(8206720, 24), to_signed(8204046, 24), to_signed(8201352, 24), to_signed(8198638, 24), to_signed(8195906, 24), to_signed(8193154, 24), to_signed(8190382, 24), to_signed(8187592, 24), to_signed(8184782, 24), to_signed(8181953, 24), to_signed(8179105, 24), to_signed(8176237, 24), to_signed(8173351, 24), to_signed(8170445, 24), to_signed(8167519, 24), to_signed(8164575, 24), to_signed(8161611, 24), to_signed(8158629, 24), to_signed(8155626, 24), to_signed(8152605, 24), to_signed(8149565, 24), to_signed(8146505, 24), to_signed(8143426, 24), to_signed(8140329, 24), to_signed(8137211, 24), to_signed(8134075, 24), to_signed(8130920, 24), to_signed(8127745, 24), to_signed(8124552, 24), to_signed(8121339, 24), to_signed(8118107, 24), to_signed(8114856, 24), to_signed(8111586, 24), to_signed(8108297, 24), to_signed(8104989, 24), to_signed(8101661, 24), to_signed(8098315, 24), to_signed(8094950, 24), to_signed(8091565, 24), to_signed(8088162, 24), to_signed(8084739, 24), to_signed(8081298, 24), to_signed(8077837, 24), to_signed(8074357, 24), to_signed(8070859, 24), to_signed(8067341, 24), to_signed(8063805, 24), to_signed(8060249, 24), to_signed(8056675, 24), to_signed(8053081, 24), to_signed(8049469, 24), to_signed(8045837, 24), to_signed(8042187, 24), to_signed(8038518, 24), to_signed(8034830, 24), to_signed(8031123, 24), to_signed(8027397, 24), to_signed(8023652, 24), to_signed(8019888, 24), to_signed(8016106, 24), to_signed(8012304, 24), to_signed(8008484, 24), to_signed(8004645, 24), to_signed(8000787, 24), to_signed(7996910, 24), to_signed(7993015, 24), to_signed(7989100, 24), to_signed(7985167, 24), to_signed(7981215, 24), to_signed(7977244, 24), to_signed(7973255, 24), to_signed(7969246, 24), to_signed(7965219, 24), to_signed(7961173, 24), to_signed(7957109, 24), to_signed(7953026, 24), to_signed(7948924, 24), to_signed(7944803, 24), to_signed(7940663, 24), to_signed(7936505, 24), to_signed(7932329, 24), to_signed(7928133, 24), to_signed(7923919, 24), to_signed(7919686, 24), to_signed(7915435, 24), to_signed(7911165, 24), to_signed(7906877, 24), to_signed(7902569, 24), to_signed(7898244, 24), to_signed(7893899, 24), to_signed(7889536, 24), to_signed(7885155, 24), to_signed(7880755, 24), to_signed(7876336, 24), to_signed(7871899, 24), to_signed(7867443, 24), to_signed(7862969, 24), to_signed(7858476, 24), to_signed(7853965, 24), to_signed(7849436, 24), to_signed(7844887, 24), to_signed(7840321, 24), to_signed(7835736, 24), to_signed(7831132, 24), to_signed(7826510, 24), to_signed(7821870, 24), to_signed(7817211, 24), to_signed(7812534, 24), to_signed(7807839, 24), to_signed(7803125, 24), to_signed(7798393, 24), to_signed(7793642, 24), to_signed(7788873, 24), to_signed(7784086, 24), to_signed(7779280, 24), to_signed(7774456, 24), to_signed(7769614, 24), to_signed(7764754, 24), to_signed(7759875, 24), to_signed(7754978, 24), to_signed(7750063, 24), to_signed(7745129, 24), to_signed(7740178, 24), to_signed(7735208, 24), to_signed(7730220, 24), to_signed(7725213, 24), to_signed(7720189, 24), to_signed(7715146, 24), to_signed(7710085, 24), to_signed(7705006, 24), to_signed(7699909, 24), to_signed(7694794, 24), to_signed(7689661, 24), to_signed(7684509, 24), to_signed(7679340, 24), to_signed(7674152, 24), to_signed(7668947, 24), to_signed(7663723, 24), to_signed(7658481, 24), to_signed(7653222, 24), to_signed(7647944, 24), to_signed(7642648, 24), to_signed(7637335, 24), to_signed(7632003, 24), to_signed(7626653, 24), to_signed(7621286, 24), to_signed(7615900, 24), to_signed(7610497, 24), to_signed(7605075, 24), to_signed(7599636, 24), to_signed(7594179, 24), to_signed(7588704, 24), to_signed(7583211, 24), to_signed(7577701, 24), to_signed(7572172, 24), to_signed(7566626, 24), to_signed(7561062, 24), to_signed(7555480, 24), to_signed(7549880, 24), to_signed(7544263, 24), to_signed(7538627, 24), to_signed(7532974, 24), to_signed(7527304, 24), to_signed(7521615, 24), to_signed(7515909, 24), to_signed(7510185, 24), to_signed(7504444, 24), to_signed(7498685, 24), to_signed(7492908, 24), to_signed(7487114, 24), to_signed(7481302, 24), to_signed(7475472, 24), to_signed(7469625, 24), to_signed(7463760, 24), to_signed(7457878, 24), to_signed(7451978, 24), to_signed(7446060, 24), to_signed(7440125, 24), to_signed(7434173, 24), to_signed(7428203, 24), to_signed(7422216, 24), to_signed(7416211, 24), to_signed(7410188, 24), to_signed(7404148, 24), to_signed(7398091, 24), to_signed(7392017, 24), to_signed(7385925, 24), to_signed(7379815, 24), to_signed(7373688, 24), to_signed(7367544, 24), to_signed(7361383, 24), to_signed(7355204, 24), to_signed(7349008, 24), to_signed(7342795, 24), to_signed(7336564, 24), to_signed(7330316, 24), to_signed(7324051, 24), to_signed(7317769, 24), to_signed(7311469, 24), to_signed(7305152, 24), to_signed(7298818, 24), to_signed(7292467, 24), to_signed(7286099, 24), to_signed(7279713, 24), to_signed(7273311, 24), to_signed(7266891, 24), to_signed(7260454, 24), to_signed(7254000, 24), to_signed(7247529, 24), to_signed(7241041, 24), to_signed(7234536, 24), to_signed(7228014, 24), to_signed(7221475, 24), to_signed(7214919, 24), to_signed(7208346, 24), to_signed(7201756, 24), to_signed(7195149, 24), to_signed(7188525, 24), to_signed(7181884, 24), to_signed(7175226, 24), to_signed(7168551, 24), to_signed(7161860, 24), to_signed(7155152, 24), to_signed(7148426, 24), to_signed(7141684, 24), to_signed(7134926, 24), to_signed(7128150, 24), to_signed(7121358, 24), to_signed(7114549, 24), to_signed(7107723, 24), to_signed(7100880, 24), to_signed(7094021, 24), to_signed(7087145, 24), to_signed(7080252, 24), to_signed(7073343, 24), to_signed(7066417, 24), to_signed(7059474, 24), to_signed(7052515, 24), to_signed(7045539, 24), to_signed(7038547, 24), to_signed(7031538, 24), to_signed(7024512, 24), to_signed(7017470, 24), to_signed(7010412, 24), to_signed(7003337, 24), to_signed(6996245, 24), to_signed(6989137, 24), to_signed(6982013, 24), to_signed(6974872, 24), to_signed(6967715, 24), to_signed(6960541, 24), to_signed(6953351, 24), to_signed(6946145, 24), to_signed(6938922, 24), to_signed(6931683, 24), to_signed(6924428, 24), to_signed(6917156, 24), to_signed(6909868, 24), to_signed(6902564, 24), to_signed(6895243, 24), to_signed(6887907, 24), to_signed(6880554, 24), to_signed(6873185, 24), to_signed(6865799, 24), to_signed(6858398, 24), to_signed(6850980, 24), to_signed(6843547, 24), to_signed(6836097, 24), to_signed(6828631, 24), to_signed(6821149, 24), to_signed(6813651, 24), to_signed(6806137, 24), to_signed(6798607, 24), to_signed(6791061, 24), to_signed(6783499, 24), to_signed(6775921, 24), to_signed(6768327, 24), to_signed(6760718, 24), to_signed(6753092, 24), to_signed(6745450, 24), to_signed(6737793, 24), to_signed(6730119, 24), to_signed(6722430, 24), to_signed(6714725, 24), to_signed(6707004, 24), to_signed(6699268, 24), to_signed(6691515, 24), to_signed(6683747, 24), to_signed(6675963, 24), to_signed(6668164, 24), to_signed(6660349, 24), to_signed(6652518, 24), to_signed(6644671, 24), to_signed(6636809, 24), to_signed(6628931, 24), to_signed(6621038, 24), to_signed(6613129, 24), to_signed(6605204, 24), to_signed(6597264, 24), to_signed(6589308, 24), to_signed(6581337, 24), to_signed(6573351, 24), to_signed(6565349, 24), to_signed(6557331, 24), to_signed(6549298, 24), to_signed(6541250, 24), to_signed(6533186, 24), to_signed(6525107, 24), to_signed(6517012, 24), to_signed(6508902, 24), to_signed(6500777, 24), to_signed(6492637, 24), to_signed(6484481, 24), to_signed(6476310, 24), to_signed(6468124, 24), to_signed(6459923, 24), to_signed(6451706, 24), to_signed(6443474, 24), to_signed(6435227, 24), to_signed(6426965, 24), to_signed(6418688, 24), to_signed(6410395, 24), to_signed(6402088, 24), to_signed(6393765, 24), to_signed(6385428, 24), to_signed(6377075, 24), to_signed(6368708, 24), to_signed(6360325, 24), to_signed(6351928, 24), to_signed(6343515, 24), to_signed(6335088, 24), to_signed(6326646, 24), to_signed(6318188, 24), to_signed(6309716, 24), to_signed(6301229, 24), to_signed(6292728, 24), to_signed(6284211, 24), to_signed(6275680, 24), to_signed(6267134, 24), to_signed(6258573, 24), to_signed(6249997, 24), to_signed(6241407, 24), to_signed(6232802, 24), to_signed(6224182, 24), to_signed(6215548, 24), to_signed(6206899, 24), to_signed(6198236, 24), to_signed(6189558, 24), to_signed(6180865, 24), to_signed(6172158, 24), to_signed(6163436, 24), to_signed(6154700, 24), to_signed(6145949, 24), to_signed(6137184, 24), to_signed(6128404, 24), to_signed(6119610, 24), to_signed(6110802, 24), to_signed(6101979, 24), to_signed(6093142, 24), to_signed(6084290, 24), to_signed(6075424, 24), to_signed(6066544, 24), to_signed(6057650, 24), to_signed(6048741, 24), to_signed(6039818, 24), to_signed(6030881, 24), to_signed(6021930, 24), to_signed(6012964, 24), to_signed(6003985, 24), to_signed(5994991, 24), to_signed(5985983, 24), to_signed(5976961, 24), to_signed(5967925, 24), to_signed(5958875, 24), to_signed(5949811, 24), to_signed(5940733, 24), to_signed(5931641, 24), to_signed(5922535, 24), to_signed(5913415, 24), to_signed(5904281, 24), to_signed(5895134, 24), to_signed(5885972, 24), to_signed(5876796, 24), to_signed(5867607, 24), to_signed(5858404, 24), to_signed(5849187, 24), to_signed(5839957, 24), to_signed(5830712, 24), to_signed(5821454, 24), to_signed(5812182, 24), to_signed(5802897, 24), to_signed(5793598, 24), to_signed(5784285, 24), to_signed(5774958, 24), to_signed(5765618, 24), to_signed(5756265, 24), to_signed(5746898, 24), to_signed(5737517, 24), to_signed(5728123, 24), to_signed(5718716, 24), to_signed(5709294, 24), to_signed(5699860, 24), to_signed(5690412, 24), to_signed(5680951, 24), to_signed(5671476, 24), to_signed(5661988, 24), to_signed(5652487, 24), to_signed(5642972, 24), to_signed(5633444, 24), to_signed(5623903, 24), to_signed(5614349, 24), to_signed(5604781, 24), to_signed(5595200, 24), to_signed(5585606, 24), to_signed(5575999, 24), to_signed(5566379, 24), to_signed(5556746, 24), to_signed(5547099, 24), to_signed(5537440, 24), to_signed(5527767, 24), to_signed(5518082, 24), to_signed(5508384, 24), to_signed(5498672, 24), to_signed(5488948, 24), to_signed(5479210, 24), to_signed(5469460, 24), to_signed(5459697, 24), to_signed(5449921, 24), to_signed(5440133, 24), to_signed(5430331, 24), to_signed(5420517, 24), to_signed(5410690, 24), to_signed(5400850, 24), to_signed(5390997, 24), to_signed(5381132, 24), to_signed(5371254, 24), to_signed(5361364, 24), to_signed(5351461, 24), to_signed(5341545, 24), to_signed(5331617, 24), to_signed(5321676, 24), to_signed(5311723, 24), to_signed(5301757, 24), to_signed(5291779, 24), to_signed(5281788, 24), to_signed(5271785, 24), to_signed(5261769, 24), to_signed(5251741, 24), to_signed(5241701, 24), to_signed(5231648, 24), to_signed(5221583, 24), to_signed(5211506, 24), to_signed(5201416, 24), to_signed(5191315, 24), to_signed(5181201, 24), to_signed(5171074, 24), to_signed(5160936, 24), to_signed(5150786, 24), to_signed(5140623, 24), to_signed(5130448, 24), to_signed(5120262, 24), to_signed(5110063, 24), to_signed(5099852, 24), to_signed(5089629, 24), to_signed(5079394, 24), to_signed(5069147, 24), to_signed(5058889, 24), to_signed(5048618, 24), to_signed(5038336, 24), to_signed(5028041, 24), to_signed(5017735, 24), to_signed(5007417, 24), to_signed(4997087, 24), to_signed(4986746, 24), to_signed(4976393, 24), to_signed(4966028, 24), to_signed(4955651, 24), to_signed(4945263, 24), to_signed(4934863, 24), to_signed(4924451, 24), to_signed(4914028, 24), to_signed(4903593, 24), to_signed(4893147, 24), to_signed(4882689, 24), to_signed(4872220, 24), to_signed(4861739, 24), to_signed(4851247, 24), to_signed(4840744, 24), to_signed(4830229, 24), to_signed(4819702, 24), to_signed(4809165, 24), to_signed(4798616, 24), to_signed(4788055, 24), to_signed(4777484, 24), to_signed(4766901, 24), to_signed(4756307, 24), to_signed(4745702, 24), to_signed(4735086, 24), to_signed(4724458, 24), to_signed(4713819, 24), to_signed(4703170, 24), to_signed(4692509, 24), to_signed(4681837, 24), to_signed(4671154, 24), to_signed(4660460, 24), to_signed(4649756, 24), to_signed(4639040, 24), to_signed(4628313, 24), to_signed(4617576, 24), to_signed(4606827, 24), to_signed(4596068, 24), to_signed(4585298, 24), to_signed(4574517, 24), to_signed(4563725, 24), to_signed(4552923, 24), to_signed(4542110, 24), to_signed(4531286, 24), to_signed(4520452, 24), to_signed(4509607, 24), to_signed(4498751, 24), to_signed(4487885, 24), to_signed(4477008, 24), to_signed(4466121, 24), to_signed(4455223, 24), to_signed(4444314, 24), to_signed(4433396, 24), to_signed(4422466, 24), to_signed(4411527, 24), to_signed(4400577, 24), to_signed(4389616, 24), to_signed(4378646, 24), to_signed(4367665, 24), to_signed(4356673, 24), to_signed(4345672, 24), to_signed(4334660, 24), to_signed(4323638, 24), to_signed(4312606, 24), to_signed(4301564, 24), to_signed(4290511, 24), to_signed(4279449, 24), to_signed(4268376, 24), to_signed(4257293, 24), to_signed(4246201, 24), to_signed(4235098, 24), to_signed(4223986, 24), to_signed(4212863, 24), to_signed(4201731, 24), to_signed(4190588, 24), to_signed(4179436, 24), to_signed(4168274, 24), to_signed(4157102, 24), to_signed(4145921, 24), to_signed(4134729, 24), to_signed(4123528, 24), to_signed(4112317, 24), to_signed(4101097, 24), to_signed(4089867, 24), to_signed(4078627, 24), to_signed(4067378, 24), to_signed(4056119, 24), to_signed(4044850, 24), to_signed(4033572, 24), to_signed(4022285, 24), to_signed(4010988, 24), to_signed(3999681, 24), to_signed(3988366, 24), to_signed(3977040, 24), to_signed(3965706, 24), to_signed(3954362, 24), to_signed(3943009, 24), to_signed(3931646, 24), to_signed(3920275, 24), to_signed(3908894, 24), to_signed(3897504, 24), to_signed(3886104, 24), to_signed(3874696, 24), to_signed(3863278, 24), to_signed(3851852, 24), to_signed(3840416, 24), to_signed(3828971, 24), to_signed(3817517, 24), to_signed(3806055, 24), to_signed(3794583, 24), to_signed(3783102, 24), to_signed(3771613, 24), to_signed(3760114, 24), to_signed(3748607, 24), to_signed(3737091, 24), to_signed(3725566, 24), to_signed(3714032, 24), to_signed(3702490, 24), to_signed(3690939, 24), to_signed(3679379, 24), to_signed(3667811, 24), to_signed(3656234, 24), to_signed(3644648, 24), to_signed(3633054, 24), to_signed(3621451, 24), to_signed(3609840, 24), to_signed(3598220, 24), to_signed(3586592, 24), to_signed(3574955, 24), to_signed(3563310, 24), to_signed(3551656, 24), to_signed(3539994, 24), to_signed(3528324, 24), to_signed(3516646, 24), to_signed(3504959, 24), to_signed(3493264, 24), to_signed(3481561, 24), to_signed(3469849, 24), to_signed(3458130, 24), to_signed(3446402, 24), to_signed(3434666, 24), to_signed(3422922, 24), to_signed(3411170, 24), to_signed(3399410, 24), to_signed(3387642, 24), to_signed(3375866, 24), to_signed(3364082, 24), to_signed(3352290, 24), to_signed(3340491, 24), to_signed(3328683, 24), to_signed(3316868, 24), to_signed(3305044, 24), to_signed(3293213, 24), to_signed(3281375, 24), to_signed(3269528, 24), to_signed(3257674, 24), to_signed(3245812, 24), to_signed(3233943, 24), to_signed(3222065, 24), to_signed(3210181, 24), to_signed(3198289, 24), to_signed(3186389, 24), to_signed(3174482, 24), to_signed(3162567, 24), to_signed(3150645, 24), to_signed(3138715, 24), to_signed(3126778, 24), to_signed(3114834, 24), to_signed(3102882, 24), to_signed(3090923, 24), to_signed(3078957, 24), to_signed(3066984, 24), to_signed(3055003, 24), to_signed(3043015, 24), to_signed(3031020, 24), to_signed(3019018, 24), to_signed(3007009, 24), to_signed(2994992, 24), to_signed(2982969, 24), to_signed(2970938, 24), to_signed(2958901, 24), to_signed(2946857, 24), to_signed(2934805, 24), to_signed(2922747, 24), to_signed(2910682, 24), to_signed(2898610, 24), to_signed(2886531, 24), to_signed(2874446, 24), to_signed(2862354, 24), to_signed(2850255, 24), to_signed(2838149, 24), to_signed(2826036, 24), to_signed(2813917, 24), to_signed(2801792, 24), to_signed(2789659, 24), to_signed(2777521, 24), to_signed(2765375, 24), to_signed(2753223, 24), to_signed(2741065, 24), to_signed(2728900, 24), to_signed(2716729, 24), to_signed(2704551, 24), to_signed(2692367, 24), to_signed(2680177, 24), to_signed(2667980, 24), to_signed(2655777, 24), to_signed(2643568, 24), to_signed(2631353, 24), to_signed(2619131, 24), to_signed(2606903, 24), to_signed(2594669, 24), to_signed(2582429, 24), to_signed(2570183, 24), to_signed(2557931, 24), to_signed(2545673, 24), to_signed(2533409, 24), to_signed(2521139, 24), to_signed(2508863, 24), to_signed(2496581, 24), to_signed(2484293, 24), to_signed(2472000, 24), to_signed(2459700, 24), to_signed(2447395, 24), to_signed(2435084, 24), to_signed(2422767, 24), to_signed(2410445, 24), to_signed(2398117, 24), to_signed(2385783, 24), to_signed(2373443, 24), to_signed(2361099, 24), to_signed(2348748, 24), to_signed(2336392, 24), to_signed(2324030, 24), to_signed(2311663, 24), to_signed(2299291, 24), to_signed(2286913, 24), to_signed(2274530, 24), to_signed(2262141, 24), to_signed(2249747, 24), to_signed(2237348, 24), to_signed(2224944, 24), to_signed(2212534, 24), to_signed(2200119, 24), to_signed(2187699, 24), to_signed(2175274, 24), to_signed(2162844, 24), to_signed(2150408, 24), to_signed(2137968, 24), to_signed(2125522, 24), to_signed(2113072, 24), to_signed(2100616, 24), to_signed(2088156, 24), to_signed(2075690, 24), to_signed(2063220, 24), to_signed(2050745, 24), to_signed(2038265, 24), to_signed(2025780, 24), to_signed(2013291, 24), to_signed(2000797, 24), to_signed(1988298, 24), to_signed(1975794, 24), to_signed(1963286, 24), to_signed(1950773, 24), to_signed(1938255, 24), to_signed(1925733, 24), to_signed(1913207, 24), to_signed(1900676, 24), to_signed(1888140, 24), to_signed(1875600, 24), to_signed(1863056, 24), to_signed(1850507, 24), to_signed(1837954, 24), to_signed(1825396, 24), to_signed(1812835, 24), to_signed(1800269, 24), to_signed(1787698, 24), to_signed(1775124, 24), to_signed(1762545, 24), to_signed(1749963, 24), to_signed(1737376, 24), to_signed(1724785, 24), to_signed(1712190, 24), to_signed(1699591, 24), to_signed(1686987, 24), to_signed(1674380, 24), to_signed(1661769, 24), to_signed(1649155, 24), to_signed(1636536, 24), to_signed(1623913, 24), to_signed(1611287, 24), to_signed(1598656, 24), to_signed(1586022, 24), to_signed(1573385, 24), to_signed(1560743, 24), to_signed(1548098, 24), to_signed(1535449, 24), to_signed(1522797, 24), to_signed(1510141, 24), to_signed(1497482, 24), to_signed(1484819, 24), to_signed(1472152, 24), to_signed(1459482, 24), to_signed(1446809, 24), to_signed(1434132, 24), to_signed(1421452, 24), to_signed(1408768, 24), to_signed(1396081, 24), to_signed(1383391, 24), to_signed(1370698, 24), to_signed(1358001, 24), to_signed(1345301, 24), to_signed(1332598, 24), to_signed(1319892, 24), to_signed(1307183, 24), to_signed(1294471, 24), to_signed(1281755, 24), to_signed(1269037, 24), to_signed(1256315, 24), to_signed(1243591, 24), to_signed(1230864, 24), to_signed(1218134, 24), to_signed(1205401, 24), to_signed(1192665, 24), to_signed(1179926, 24), to_signed(1167185, 24), to_signed(1154441, 24), to_signed(1141694, 24), to_signed(1128944, 24), to_signed(1116192, 24), to_signed(1103437, 24), to_signed(1090680, 24), to_signed(1077920, 24), to_signed(1065157, 24), to_signed(1052392, 24), to_signed(1039625, 24), to_signed(1026855, 24), to_signed(1014082, 24), to_signed(1001307, 24), to_signed(988530, 24), to_signed(975751, 24), to_signed(962969, 24), to_signed(950185, 24), to_signed(937399, 24), to_signed(924610, 24), to_signed(911820, 24), to_signed(899027, 24), to_signed(886232, 24), to_signed(873435, 24), to_signed(860636, 24), to_signed(847835, 24), to_signed(835032, 24), to_signed(822227, 24), to_signed(809420, 24), to_signed(796611, 24), to_signed(783800, 24), to_signed(770988, 24), to_signed(758173, 24), to_signed(745357, 24), to_signed(732539, 24), to_signed(719720, 24), to_signed(706898, 24), to_signed(694075, 24), to_signed(681250, 24), to_signed(668424, 24), to_signed(655596, 24), to_signed(642767, 24), to_signed(629936, 24), to_signed(617104, 24), to_signed(604270, 24), to_signed(591435, 24), to_signed(578598, 24), to_signed(565760, 24), to_signed(552921, 24), to_signed(540080, 24), to_signed(527238, 24), to_signed(514395, 24), to_signed(501551, 24), to_signed(488705, 24), to_signed(475859, 24), to_signed(463011, 24), to_signed(450162, 24), to_signed(437312, 24), to_signed(424461, 24), to_signed(411609, 24), to_signed(398756, 24), to_signed(385902, 24), to_signed(373047, 24), to_signed(360192, 24), to_signed(347335, 24), to_signed(334478, 24), to_signed(321620, 24), to_signed(308761, 24), to_signed(295901, 24), to_signed(283041, 24), to_signed(270180, 24), to_signed(257318, 24), to_signed(244456, 24), to_signed(231593, 24), to_signed(218730, 24), to_signed(205866, 24), to_signed(193002, 24), to_signed(180137, 24), to_signed(167272, 24), to_signed(154406, 24), to_signed(141540, 24), to_signed(128674, 24), to_signed(115807, 24), to_signed(102941, 24), to_signed(90074, 24), to_signed(77206, 24), to_signed(64339, 24), to_signed(51471, 24), to_signed(38603, 24), to_signed(25735, 24), to_signed(12867, 24), to_signed(0, 24), to_signed(-12867, 24), to_signed(-25735, 24), to_signed(-38603, 24), to_signed(-51471, 24), to_signed(-64339, 24), to_signed(-77206, 24), to_signed(-90074, 24), to_signed(-102941, 24), to_signed(-115807, 24), to_signed(-128674, 24), to_signed(-141540, 24), to_signed(-154406, 24), to_signed(-167272, 24), to_signed(-180137, 24), to_signed(-193002, 24), to_signed(-205866, 24), to_signed(-218730, 24), to_signed(-231593, 24), to_signed(-244456, 24), to_signed(-257318, 24), to_signed(-270180, 24), to_signed(-283041, 24), to_signed(-295901, 24), to_signed(-308761, 24), to_signed(-321620, 24), to_signed(-334478, 24), to_signed(-347335, 24), to_signed(-360192, 24), to_signed(-373047, 24), to_signed(-385902, 24), to_signed(-398756, 24), to_signed(-411609, 24), to_signed(-424461, 24), to_signed(-437312, 24), to_signed(-450162, 24), to_signed(-463011, 24), to_signed(-475859, 24), to_signed(-488705, 24), to_signed(-501551, 24), to_signed(-514395, 24), to_signed(-527238, 24), to_signed(-540080, 24), to_signed(-552921, 24), to_signed(-565760, 24), to_signed(-578598, 24), to_signed(-591435, 24), to_signed(-604270, 24), to_signed(-617104, 24), to_signed(-629936, 24), to_signed(-642767, 24), to_signed(-655596, 24), to_signed(-668424, 24), to_signed(-681250, 24), to_signed(-694075, 24), to_signed(-706898, 24), to_signed(-719720, 24), to_signed(-732539, 24), to_signed(-745357, 24), to_signed(-758173, 24), to_signed(-770988, 24), to_signed(-783800, 24), to_signed(-796611, 24), to_signed(-809420, 24), to_signed(-822227, 24), to_signed(-835032, 24), to_signed(-847835, 24), to_signed(-860636, 24), to_signed(-873435, 24), to_signed(-886232, 24), to_signed(-899027, 24), to_signed(-911820, 24), to_signed(-924610, 24), to_signed(-937399, 24), to_signed(-950185, 24), to_signed(-962969, 24), to_signed(-975751, 24), to_signed(-988530, 24), to_signed(-1001307, 24), to_signed(-1014082, 24), to_signed(-1026855, 24), to_signed(-1039625, 24), to_signed(-1052392, 24), to_signed(-1065157, 24), to_signed(-1077920, 24), to_signed(-1090680, 24), to_signed(-1103437, 24), to_signed(-1116192, 24), to_signed(-1128944, 24), to_signed(-1141694, 24), to_signed(-1154441, 24), to_signed(-1167185, 24), to_signed(-1179926, 24), to_signed(-1192665, 24), to_signed(-1205401, 24), to_signed(-1218134, 24), to_signed(-1230864, 24), to_signed(-1243591, 24), to_signed(-1256315, 24), to_signed(-1269037, 24), to_signed(-1281755, 24), to_signed(-1294471, 24), to_signed(-1307183, 24), to_signed(-1319892, 24), to_signed(-1332598, 24), to_signed(-1345301, 24), to_signed(-1358001, 24), to_signed(-1370698, 24), to_signed(-1383391, 24), to_signed(-1396081, 24), to_signed(-1408768, 24), to_signed(-1421452, 24), to_signed(-1434132, 24), to_signed(-1446809, 24), to_signed(-1459482, 24), to_signed(-1472152, 24), to_signed(-1484819, 24), to_signed(-1497482, 24), to_signed(-1510141, 24), to_signed(-1522797, 24), to_signed(-1535449, 24), to_signed(-1548098, 24), to_signed(-1560743, 24), to_signed(-1573385, 24), to_signed(-1586022, 24), to_signed(-1598656, 24), to_signed(-1611287, 24), to_signed(-1623913, 24), to_signed(-1636536, 24), to_signed(-1649155, 24), to_signed(-1661769, 24), to_signed(-1674380, 24), to_signed(-1686987, 24), to_signed(-1699591, 24), to_signed(-1712190, 24), to_signed(-1724785, 24), to_signed(-1737376, 24), to_signed(-1749963, 24), to_signed(-1762545, 24), to_signed(-1775124, 24), to_signed(-1787698, 24), to_signed(-1800269, 24), to_signed(-1812835, 24), to_signed(-1825396, 24), to_signed(-1837954, 24), to_signed(-1850507, 24), to_signed(-1863056, 24), to_signed(-1875600, 24), to_signed(-1888140, 24), to_signed(-1900676, 24), to_signed(-1913207, 24), to_signed(-1925733, 24), to_signed(-1938255, 24), to_signed(-1950773, 24), to_signed(-1963286, 24), to_signed(-1975794, 24), to_signed(-1988298, 24), to_signed(-2000797, 24), to_signed(-2013291, 24), to_signed(-2025780, 24), to_signed(-2038265, 24), to_signed(-2050745, 24), to_signed(-2063220, 24), to_signed(-2075690, 24), to_signed(-2088156, 24), to_signed(-2100616, 24), to_signed(-2113072, 24), to_signed(-2125522, 24), to_signed(-2137968, 24), to_signed(-2150408, 24), to_signed(-2162844, 24), to_signed(-2175274, 24), to_signed(-2187699, 24), to_signed(-2200119, 24), to_signed(-2212534, 24), to_signed(-2224944, 24), to_signed(-2237348, 24), to_signed(-2249747, 24), to_signed(-2262141, 24), to_signed(-2274530, 24), to_signed(-2286913, 24), to_signed(-2299291, 24), to_signed(-2311663, 24), to_signed(-2324030, 24), to_signed(-2336392, 24), to_signed(-2348748, 24), to_signed(-2361099, 24), to_signed(-2373443, 24), to_signed(-2385783, 24), to_signed(-2398117, 24), to_signed(-2410445, 24), to_signed(-2422767, 24), to_signed(-2435084, 24), to_signed(-2447395, 24), to_signed(-2459700, 24), to_signed(-2472000, 24), to_signed(-2484293, 24), to_signed(-2496581, 24), to_signed(-2508863, 24), to_signed(-2521139, 24), to_signed(-2533409, 24), to_signed(-2545673, 24), to_signed(-2557931, 24), to_signed(-2570183, 24), to_signed(-2582429, 24), to_signed(-2594669, 24), to_signed(-2606903, 24), to_signed(-2619131, 24), to_signed(-2631353, 24), to_signed(-2643568, 24), to_signed(-2655777, 24), to_signed(-2667980, 24), to_signed(-2680177, 24), to_signed(-2692367, 24), to_signed(-2704551, 24), to_signed(-2716729, 24), to_signed(-2728900, 24), to_signed(-2741065, 24), to_signed(-2753223, 24), to_signed(-2765375, 24), to_signed(-2777521, 24), to_signed(-2789659, 24), to_signed(-2801792, 24), to_signed(-2813917, 24), to_signed(-2826036, 24), to_signed(-2838149, 24), to_signed(-2850255, 24), to_signed(-2862354, 24), to_signed(-2874446, 24), to_signed(-2886531, 24), to_signed(-2898610, 24), to_signed(-2910682, 24), to_signed(-2922747, 24), to_signed(-2934805, 24), to_signed(-2946857, 24), to_signed(-2958901, 24), to_signed(-2970938, 24), to_signed(-2982969, 24), to_signed(-2994992, 24), to_signed(-3007009, 24), to_signed(-3019018, 24), to_signed(-3031020, 24), to_signed(-3043015, 24), to_signed(-3055003, 24), to_signed(-3066984, 24), to_signed(-3078957, 24), to_signed(-3090923, 24), to_signed(-3102882, 24), to_signed(-3114834, 24), to_signed(-3126778, 24), to_signed(-3138715, 24), to_signed(-3150645, 24), to_signed(-3162567, 24), to_signed(-3174482, 24), to_signed(-3186389, 24), to_signed(-3198289, 24), to_signed(-3210181, 24), to_signed(-3222065, 24), to_signed(-3233943, 24), to_signed(-3245812, 24), to_signed(-3257674, 24), to_signed(-3269528, 24), to_signed(-3281375, 24), to_signed(-3293213, 24), to_signed(-3305044, 24), to_signed(-3316868, 24), to_signed(-3328683, 24), to_signed(-3340491, 24), to_signed(-3352290, 24), to_signed(-3364082, 24), to_signed(-3375866, 24), to_signed(-3387642, 24), to_signed(-3399410, 24), to_signed(-3411170, 24), to_signed(-3422922, 24), to_signed(-3434666, 24), to_signed(-3446402, 24), to_signed(-3458130, 24), to_signed(-3469849, 24), to_signed(-3481561, 24), to_signed(-3493264, 24), to_signed(-3504959, 24), to_signed(-3516646, 24), to_signed(-3528324, 24), to_signed(-3539994, 24), to_signed(-3551656, 24), to_signed(-3563310, 24), to_signed(-3574955, 24), to_signed(-3586592, 24), to_signed(-3598220, 24), to_signed(-3609840, 24), to_signed(-3621451, 24), to_signed(-3633054, 24), to_signed(-3644648, 24), to_signed(-3656234, 24), to_signed(-3667811, 24), to_signed(-3679379, 24), to_signed(-3690939, 24), to_signed(-3702490, 24), to_signed(-3714032, 24), to_signed(-3725566, 24), to_signed(-3737091, 24), to_signed(-3748607, 24), to_signed(-3760114, 24), to_signed(-3771613, 24), to_signed(-3783102, 24), to_signed(-3794583, 24), to_signed(-3806055, 24), to_signed(-3817517, 24), to_signed(-3828971, 24), to_signed(-3840416, 24), to_signed(-3851852, 24), to_signed(-3863278, 24), to_signed(-3874696, 24), to_signed(-3886104, 24), to_signed(-3897504, 24), to_signed(-3908894, 24), to_signed(-3920275, 24), to_signed(-3931646, 24), to_signed(-3943009, 24), to_signed(-3954362, 24), to_signed(-3965706, 24), to_signed(-3977040, 24), to_signed(-3988366, 24), to_signed(-3999681, 24), to_signed(-4010988, 24), to_signed(-4022285, 24), to_signed(-4033572, 24), to_signed(-4044850, 24), to_signed(-4056119, 24), to_signed(-4067378, 24), to_signed(-4078627, 24), to_signed(-4089867, 24), to_signed(-4101097, 24), to_signed(-4112317, 24), to_signed(-4123528, 24), to_signed(-4134729, 24), to_signed(-4145921, 24), to_signed(-4157102, 24), to_signed(-4168274, 24), to_signed(-4179436, 24), to_signed(-4190588, 24), to_signed(-4201731, 24), to_signed(-4212863, 24), to_signed(-4223986, 24), to_signed(-4235098, 24), to_signed(-4246201, 24), to_signed(-4257293, 24), to_signed(-4268376, 24), to_signed(-4279449, 24), to_signed(-4290511, 24), to_signed(-4301564, 24), to_signed(-4312606, 24), to_signed(-4323638, 24), to_signed(-4334660, 24), to_signed(-4345672, 24), to_signed(-4356673, 24), to_signed(-4367665, 24), to_signed(-4378646, 24), to_signed(-4389616, 24), to_signed(-4400577, 24), to_signed(-4411527, 24), to_signed(-4422466, 24), to_signed(-4433396, 24), to_signed(-4444314, 24), to_signed(-4455223, 24), to_signed(-4466121, 24), to_signed(-4477008, 24), to_signed(-4487885, 24), to_signed(-4498751, 24), to_signed(-4509607, 24), to_signed(-4520452, 24), to_signed(-4531286, 24), to_signed(-4542110, 24), to_signed(-4552923, 24), to_signed(-4563725, 24), to_signed(-4574517, 24), to_signed(-4585298, 24), to_signed(-4596068, 24), to_signed(-4606827, 24), to_signed(-4617576, 24), to_signed(-4628313, 24), to_signed(-4639040, 24), to_signed(-4649756, 24), to_signed(-4660460, 24), to_signed(-4671154, 24), to_signed(-4681837, 24), to_signed(-4692509, 24), to_signed(-4703170, 24), to_signed(-4713819, 24), to_signed(-4724458, 24), to_signed(-4735086, 24), to_signed(-4745702, 24), to_signed(-4756307, 24), to_signed(-4766901, 24), to_signed(-4777484, 24), to_signed(-4788055, 24), to_signed(-4798616, 24), to_signed(-4809165, 24), to_signed(-4819702, 24), to_signed(-4830229, 24), to_signed(-4840744, 24), to_signed(-4851247, 24), to_signed(-4861739, 24), to_signed(-4872220, 24), to_signed(-4882689, 24), to_signed(-4893147, 24), to_signed(-4903593, 24), to_signed(-4914028, 24), to_signed(-4924451, 24), to_signed(-4934863, 24), to_signed(-4945263, 24), to_signed(-4955651, 24), to_signed(-4966028, 24), to_signed(-4976393, 24), to_signed(-4986746, 24), to_signed(-4997087, 24), to_signed(-5007417, 24), to_signed(-5017735, 24), to_signed(-5028041, 24), to_signed(-5038336, 24), to_signed(-5048618, 24), to_signed(-5058889, 24), to_signed(-5069147, 24), to_signed(-5079394, 24), to_signed(-5089629, 24), to_signed(-5099852, 24), to_signed(-5110063, 24), to_signed(-5120262, 24), to_signed(-5130448, 24), to_signed(-5140623, 24), to_signed(-5150786, 24), to_signed(-5160936, 24), to_signed(-5171074, 24), to_signed(-5181201, 24), to_signed(-5191315, 24), to_signed(-5201416, 24), to_signed(-5211506, 24), to_signed(-5221583, 24), to_signed(-5231648, 24), to_signed(-5241701, 24), to_signed(-5251741, 24), to_signed(-5261769, 24), to_signed(-5271785, 24), to_signed(-5281788, 24), to_signed(-5291779, 24), to_signed(-5301757, 24), to_signed(-5311723, 24), to_signed(-5321676, 24), to_signed(-5331617, 24), to_signed(-5341545, 24), to_signed(-5351461, 24), to_signed(-5361364, 24), to_signed(-5371254, 24), to_signed(-5381132, 24), to_signed(-5390997, 24), to_signed(-5400850, 24), to_signed(-5410690, 24), to_signed(-5420517, 24), to_signed(-5430331, 24), to_signed(-5440133, 24), to_signed(-5449921, 24), to_signed(-5459697, 24), to_signed(-5469460, 24), to_signed(-5479210, 24), to_signed(-5488948, 24), to_signed(-5498672, 24), to_signed(-5508384, 24), to_signed(-5518082, 24), to_signed(-5527767, 24), to_signed(-5537440, 24), to_signed(-5547099, 24), to_signed(-5556746, 24), to_signed(-5566379, 24), to_signed(-5575999, 24), to_signed(-5585606, 24), to_signed(-5595200, 24), to_signed(-5604781, 24), to_signed(-5614349, 24), to_signed(-5623903, 24), to_signed(-5633444, 24), to_signed(-5642972, 24), to_signed(-5652487, 24), to_signed(-5661988, 24), to_signed(-5671476, 24), to_signed(-5680951, 24), to_signed(-5690412, 24), to_signed(-5699860, 24), to_signed(-5709294, 24), to_signed(-5718716, 24), to_signed(-5728123, 24), to_signed(-5737517, 24), to_signed(-5746898, 24), to_signed(-5756265, 24), to_signed(-5765618, 24), to_signed(-5774958, 24), to_signed(-5784285, 24), to_signed(-5793598, 24), to_signed(-5802897, 24), to_signed(-5812182, 24), to_signed(-5821454, 24), to_signed(-5830712, 24), to_signed(-5839957, 24), to_signed(-5849187, 24), to_signed(-5858404, 24), to_signed(-5867607, 24), to_signed(-5876796, 24), to_signed(-5885972, 24), to_signed(-5895134, 24), to_signed(-5904281, 24), to_signed(-5913415, 24), to_signed(-5922535, 24), to_signed(-5931641, 24), to_signed(-5940733, 24), to_signed(-5949811, 24), to_signed(-5958875, 24), to_signed(-5967925, 24), to_signed(-5976961, 24), to_signed(-5985983, 24), to_signed(-5994991, 24), to_signed(-6003985, 24), to_signed(-6012964, 24), to_signed(-6021930, 24), to_signed(-6030881, 24), to_signed(-6039818, 24), to_signed(-6048741, 24), to_signed(-6057650, 24), to_signed(-6066544, 24), to_signed(-6075424, 24), to_signed(-6084290, 24), to_signed(-6093142, 24), to_signed(-6101979, 24), to_signed(-6110802, 24), to_signed(-6119610, 24), to_signed(-6128404, 24), to_signed(-6137184, 24), to_signed(-6145949, 24), to_signed(-6154700, 24), to_signed(-6163436, 24), to_signed(-6172158, 24), to_signed(-6180865, 24), to_signed(-6189558, 24), to_signed(-6198236, 24), to_signed(-6206899, 24), to_signed(-6215548, 24), to_signed(-6224182, 24), to_signed(-6232802, 24), to_signed(-6241407, 24), to_signed(-6249997, 24), to_signed(-6258573, 24), to_signed(-6267134, 24), to_signed(-6275680, 24), to_signed(-6284211, 24), to_signed(-6292728, 24), to_signed(-6301229, 24), to_signed(-6309716, 24), to_signed(-6318188, 24), to_signed(-6326646, 24), to_signed(-6335088, 24), to_signed(-6343515, 24), to_signed(-6351928, 24), to_signed(-6360325, 24), to_signed(-6368708, 24), to_signed(-6377075, 24), to_signed(-6385428, 24), to_signed(-6393765, 24), to_signed(-6402088, 24), to_signed(-6410395, 24), to_signed(-6418688, 24), to_signed(-6426965, 24), to_signed(-6435227, 24), to_signed(-6443474, 24), to_signed(-6451706, 24), to_signed(-6459923, 24), to_signed(-6468124, 24), to_signed(-6476310, 24), to_signed(-6484481, 24), to_signed(-6492637, 24), to_signed(-6500777, 24), to_signed(-6508902, 24), to_signed(-6517012, 24), to_signed(-6525107, 24), to_signed(-6533186, 24), to_signed(-6541250, 24), to_signed(-6549298, 24), to_signed(-6557331, 24), to_signed(-6565349, 24), to_signed(-6573351, 24), to_signed(-6581337, 24), to_signed(-6589308, 24), to_signed(-6597264, 24), to_signed(-6605204, 24), to_signed(-6613129, 24), to_signed(-6621038, 24), to_signed(-6628931, 24), to_signed(-6636809, 24), to_signed(-6644671, 24), to_signed(-6652518, 24), to_signed(-6660349, 24), to_signed(-6668164, 24), to_signed(-6675963, 24), to_signed(-6683747, 24), to_signed(-6691515, 24), to_signed(-6699268, 24), to_signed(-6707004, 24), to_signed(-6714725, 24), to_signed(-6722430, 24), to_signed(-6730119, 24), to_signed(-6737793, 24), to_signed(-6745450, 24), to_signed(-6753092, 24), to_signed(-6760718, 24), to_signed(-6768327, 24), to_signed(-6775921, 24), to_signed(-6783499, 24), to_signed(-6791061, 24), to_signed(-6798607, 24), to_signed(-6806137, 24), to_signed(-6813651, 24), to_signed(-6821149, 24), to_signed(-6828631, 24), to_signed(-6836097, 24), to_signed(-6843547, 24), to_signed(-6850980, 24), to_signed(-6858398, 24), to_signed(-6865799, 24), to_signed(-6873185, 24), to_signed(-6880554, 24), to_signed(-6887907, 24), to_signed(-6895243, 24), to_signed(-6902564, 24), to_signed(-6909868, 24), to_signed(-6917156, 24), to_signed(-6924428, 24), to_signed(-6931683, 24), to_signed(-6938922, 24), to_signed(-6946145, 24), to_signed(-6953351, 24), to_signed(-6960541, 24), to_signed(-6967715, 24), to_signed(-6974872, 24), to_signed(-6982013, 24), to_signed(-6989137, 24), to_signed(-6996245, 24), to_signed(-7003337, 24), to_signed(-7010412, 24), to_signed(-7017470, 24), to_signed(-7024512, 24), to_signed(-7031538, 24), to_signed(-7038547, 24), to_signed(-7045539, 24), to_signed(-7052515, 24), to_signed(-7059474, 24), to_signed(-7066417, 24), to_signed(-7073343, 24), to_signed(-7080252, 24), to_signed(-7087145, 24), to_signed(-7094021, 24), to_signed(-7100880, 24), to_signed(-7107723, 24), to_signed(-7114549, 24), to_signed(-7121358, 24), to_signed(-7128150, 24), to_signed(-7134926, 24), to_signed(-7141684, 24), to_signed(-7148426, 24), to_signed(-7155152, 24), to_signed(-7161860, 24), to_signed(-7168551, 24), to_signed(-7175226, 24), to_signed(-7181884, 24), to_signed(-7188525, 24), to_signed(-7195149, 24), to_signed(-7201756, 24), to_signed(-7208346, 24), to_signed(-7214919, 24), to_signed(-7221475, 24), to_signed(-7228014, 24), to_signed(-7234536, 24), to_signed(-7241041, 24), to_signed(-7247529, 24), to_signed(-7254000, 24), to_signed(-7260454, 24), to_signed(-7266891, 24), to_signed(-7273311, 24), to_signed(-7279713, 24), to_signed(-7286099, 24), to_signed(-7292467, 24), to_signed(-7298818, 24), to_signed(-7305152, 24), to_signed(-7311469, 24), to_signed(-7317769, 24), to_signed(-7324051, 24), to_signed(-7330316, 24), to_signed(-7336564, 24), to_signed(-7342795, 24), to_signed(-7349008, 24), to_signed(-7355204, 24), to_signed(-7361383, 24), to_signed(-7367544, 24), to_signed(-7373688, 24), to_signed(-7379815, 24), to_signed(-7385925, 24), to_signed(-7392017, 24), to_signed(-7398091, 24), to_signed(-7404148, 24), to_signed(-7410188, 24), to_signed(-7416211, 24), to_signed(-7422216, 24), to_signed(-7428203, 24), to_signed(-7434173, 24), to_signed(-7440125, 24), to_signed(-7446060, 24), to_signed(-7451978, 24), to_signed(-7457878, 24), to_signed(-7463760, 24), to_signed(-7469625, 24), to_signed(-7475472, 24), to_signed(-7481302, 24), to_signed(-7487114, 24), to_signed(-7492908, 24), to_signed(-7498685, 24), to_signed(-7504444, 24), to_signed(-7510185, 24), to_signed(-7515909, 24), to_signed(-7521615, 24), to_signed(-7527304, 24), to_signed(-7532974, 24), to_signed(-7538627, 24), to_signed(-7544263, 24), to_signed(-7549880, 24), to_signed(-7555480, 24), to_signed(-7561062, 24), to_signed(-7566626, 24), to_signed(-7572172, 24), to_signed(-7577701, 24), to_signed(-7583211, 24), to_signed(-7588704, 24), to_signed(-7594179, 24), to_signed(-7599636, 24), to_signed(-7605075, 24), to_signed(-7610497, 24), to_signed(-7615900, 24), to_signed(-7621286, 24), to_signed(-7626653, 24), to_signed(-7632003, 24), to_signed(-7637335, 24), to_signed(-7642648, 24), to_signed(-7647944, 24), to_signed(-7653222, 24), to_signed(-7658481, 24), to_signed(-7663723, 24), to_signed(-7668947, 24), to_signed(-7674152, 24), to_signed(-7679340, 24), to_signed(-7684509, 24), to_signed(-7689661, 24), to_signed(-7694794, 24), to_signed(-7699909, 24), to_signed(-7705006, 24), to_signed(-7710085, 24), to_signed(-7715146, 24), to_signed(-7720189, 24), to_signed(-7725213, 24), to_signed(-7730220, 24), to_signed(-7735208, 24), to_signed(-7740178, 24), to_signed(-7745129, 24), to_signed(-7750063, 24), to_signed(-7754978, 24), to_signed(-7759875, 24), to_signed(-7764754, 24), to_signed(-7769614, 24), to_signed(-7774456, 24), to_signed(-7779280, 24), to_signed(-7784086, 24), to_signed(-7788873, 24), to_signed(-7793642, 24), to_signed(-7798393, 24), to_signed(-7803125, 24), to_signed(-7807839, 24), to_signed(-7812534, 24), to_signed(-7817211, 24), to_signed(-7821870, 24), to_signed(-7826510, 24), to_signed(-7831132, 24), to_signed(-7835736, 24), to_signed(-7840321, 24), to_signed(-7844887, 24), to_signed(-7849436, 24), to_signed(-7853965, 24), to_signed(-7858476, 24), to_signed(-7862969, 24), to_signed(-7867443, 24), to_signed(-7871899, 24), to_signed(-7876336, 24), to_signed(-7880755, 24), to_signed(-7885155, 24), to_signed(-7889536, 24), to_signed(-7893899, 24), to_signed(-7898244, 24), to_signed(-7902569, 24), to_signed(-7906877, 24), to_signed(-7911165, 24), to_signed(-7915435, 24), to_signed(-7919686, 24), to_signed(-7923919, 24), to_signed(-7928133, 24), to_signed(-7932329, 24), to_signed(-7936505, 24), to_signed(-7940663, 24), to_signed(-7944803, 24), to_signed(-7948924, 24), to_signed(-7953026, 24), to_signed(-7957109, 24), to_signed(-7961173, 24), to_signed(-7965219, 24), to_signed(-7969246, 24), to_signed(-7973255, 24), to_signed(-7977244, 24), to_signed(-7981215, 24), to_signed(-7985167, 24), to_signed(-7989100, 24), to_signed(-7993015, 24), to_signed(-7996910, 24), to_signed(-8000787, 24), to_signed(-8004645, 24), to_signed(-8008484, 24), to_signed(-8012304, 24), to_signed(-8016106, 24), to_signed(-8019888, 24), to_signed(-8023652, 24), to_signed(-8027397, 24), to_signed(-8031123, 24), to_signed(-8034830, 24), to_signed(-8038518, 24), to_signed(-8042187, 24), to_signed(-8045837, 24), to_signed(-8049469, 24), to_signed(-8053081, 24), to_signed(-8056675, 24), to_signed(-8060249, 24), to_signed(-8063805, 24), to_signed(-8067341, 24), to_signed(-8070859, 24), to_signed(-8074357, 24), to_signed(-8077837, 24), to_signed(-8081298, 24), to_signed(-8084739, 24), to_signed(-8088162, 24), to_signed(-8091565, 24), to_signed(-8094950, 24), to_signed(-8098315, 24), to_signed(-8101661, 24), to_signed(-8104989, 24), to_signed(-8108297, 24), to_signed(-8111586, 24), to_signed(-8114856, 24), to_signed(-8118107, 24), to_signed(-8121339, 24), to_signed(-8124552, 24), to_signed(-8127745, 24), to_signed(-8130920, 24), to_signed(-8134075, 24), to_signed(-8137211, 24), to_signed(-8140329, 24), to_signed(-8143426, 24), to_signed(-8146505, 24), to_signed(-8149565, 24), to_signed(-8152605, 24), to_signed(-8155626, 24), to_signed(-8158629, 24), to_signed(-8161611, 24), to_signed(-8164575, 24), to_signed(-8167519, 24), to_signed(-8170445, 24), to_signed(-8173351, 24), to_signed(-8176237, 24), to_signed(-8179105, 24), to_signed(-8181953, 24), to_signed(-8184782, 24), to_signed(-8187592, 24), to_signed(-8190382, 24), to_signed(-8193154, 24), to_signed(-8195906, 24), to_signed(-8198638, 24), to_signed(-8201352, 24), to_signed(-8204046, 24), to_signed(-8206720, 24), to_signed(-8209376, 24), to_signed(-8212012, 24), to_signed(-8214629, 24), to_signed(-8217226, 24), to_signed(-8219804, 24), to_signed(-8222363, 24), to_signed(-8224903, 24), to_signed(-8227423, 24), to_signed(-8229923, 24), to_signed(-8232405, 24), to_signed(-8234867, 24), to_signed(-8237309, 24), to_signed(-8239733, 24), to_signed(-8242137, 24), to_signed(-8244521, 24), to_signed(-8246886, 24), to_signed(-8249232, 24), to_signed(-8251558, 24), to_signed(-8253865, 24), to_signed(-8256152, 24), to_signed(-8258420, 24), to_signed(-8260669, 24), to_signed(-8262898, 24), to_signed(-8265107, 24), to_signed(-8267298, 24), to_signed(-8269468, 24), to_signed(-8271620, 24), to_signed(-8273751, 24), to_signed(-8275864, 24), to_signed(-8277957, 24), to_signed(-8280030, 24), to_signed(-8282084, 24), to_signed(-8284119, 24), to_signed(-8286133, 24), to_signed(-8288129, 24), to_signed(-8290105, 24), to_signed(-8292061, 24), to_signed(-8293998, 24), to_signed(-8295916, 24), to_signed(-8297813, 24), to_signed(-8299692, 24), to_signed(-8301551, 24), to_signed(-8303390, 24), to_signed(-8305210, 24), to_signed(-8307010, 24), to_signed(-8308791, 24), to_signed(-8310552, 24), to_signed(-8312293, 24), to_signed(-8314015, 24), to_signed(-8315718, 24), to_signed(-8317401, 24), to_signed(-8319064, 24), to_signed(-8320708, 24), to_signed(-8322332, 24), to_signed(-8323936, 24), to_signed(-8325521, 24), to_signed(-8327087, 24), to_signed(-8328632, 24), to_signed(-8330159, 24), to_signed(-8331665, 24), to_signed(-8333152, 24), to_signed(-8334620, 24), to_signed(-8336067, 24), to_signed(-8337495, 24), to_signed(-8338904, 24), to_signed(-8340293, 24), to_signed(-8341662, 24), to_signed(-8343012, 24), to_signed(-8344342, 24), to_signed(-8345652, 24), to_signed(-8346943, 24), to_signed(-8348214, 24), to_signed(-8349466, 24), to_signed(-8350697, 24), to_signed(-8351909, 24), to_signed(-8353102, 24), to_signed(-8354275, 24), to_signed(-8355428, 24), to_signed(-8356562, 24), to_signed(-8357675, 24), to_signed(-8358770, 24), to_signed(-8359844, 24), to_signed(-8360899, 24), to_signed(-8361934, 24), to_signed(-8362950, 24), to_signed(-8363946, 24), to_signed(-8364922, 24), to_signed(-8365878, 24), to_signed(-8366815, 24), to_signed(-8367732, 24), to_signed(-8368629, 24), to_signed(-8369507, 24), to_signed(-8370365, 24), to_signed(-8371204, 24), to_signed(-8372022, 24), to_signed(-8372821, 24), to_signed(-8373600, 24), to_signed(-8374360, 24), to_signed(-8375100, 24), to_signed(-8375820, 24), to_signed(-8376520, 24), to_signed(-8377201, 24), to_signed(-8377862, 24), to_signed(-8378503, 24), to_signed(-8379125, 24), to_signed(-8379726, 24), to_signed(-8380309, 24), to_signed(-8380871, 24), to_signed(-8381414, 24), to_signed(-8381937, 24), to_signed(-8382440, 24), to_signed(-8382923, 24), to_signed(-8383387, 24), to_signed(-8383831, 24), to_signed(-8384255, 24), to_signed(-8384660, 24), to_signed(-8385045, 24), to_signed(-8385410, 24), to_signed(-8385755, 24), to_signed(-8386081, 24), to_signed(-8386387, 24), to_signed(-8386673, 24), to_signed(-8386940, 24), to_signed(-8387186, 24), to_signed(-8387413, 24), to_signed(-8387621, 24), to_signed(-8387808, 24), to_signed(-8387976, 24), to_signed(-8388124, 24), to_signed(-8388252, 24), to_signed(-8388361, 24), to_signed(-8388450, 24), to_signed(-8388519, 24), to_signed(-8388568, 24), to_signed(-8388598, 24), to_signed(-8388608, 24), to_signed(-8388598, 24), to_signed(-8388568, 24), to_signed(-8388519, 24), to_signed(-8388450, 24), to_signed(-8388361, 24), to_signed(-8388252, 24), to_signed(-8388124, 24), to_signed(-8387976, 24), to_signed(-8387808, 24), to_signed(-8387621, 24), to_signed(-8387413, 24), to_signed(-8387186, 24), to_signed(-8386940, 24), to_signed(-8386673, 24), to_signed(-8386387, 24), to_signed(-8386081, 24), to_signed(-8385755, 24), to_signed(-8385410, 24), to_signed(-8385045, 24), to_signed(-8384660, 24), to_signed(-8384255, 24), to_signed(-8383831, 24), to_signed(-8383387, 24), to_signed(-8382923, 24), to_signed(-8382440, 24), to_signed(-8381937, 24), to_signed(-8381414, 24), to_signed(-8380871, 24), to_signed(-8380309, 24), to_signed(-8379726, 24), to_signed(-8379125, 24), to_signed(-8378503, 24), to_signed(-8377862, 24), to_signed(-8377201, 24), to_signed(-8376520, 24), to_signed(-8375820, 24), to_signed(-8375100, 24), to_signed(-8374360, 24), to_signed(-8373600, 24), to_signed(-8372821, 24), to_signed(-8372022, 24), to_signed(-8371204, 24), to_signed(-8370365, 24), to_signed(-8369507, 24), to_signed(-8368629, 24), to_signed(-8367732, 24), to_signed(-8366815, 24), to_signed(-8365878, 24), to_signed(-8364922, 24), to_signed(-8363946, 24), to_signed(-8362950, 24), to_signed(-8361934, 24), to_signed(-8360899, 24), to_signed(-8359844, 24), to_signed(-8358770, 24), to_signed(-8357675, 24), to_signed(-8356562, 24), to_signed(-8355428, 24), to_signed(-8354275, 24), to_signed(-8353102, 24), to_signed(-8351909, 24), to_signed(-8350697, 24), to_signed(-8349466, 24), to_signed(-8348214, 24), to_signed(-8346943, 24), to_signed(-8345652, 24), to_signed(-8344342, 24), to_signed(-8343012, 24), to_signed(-8341662, 24), to_signed(-8340293, 24), to_signed(-8338904, 24), to_signed(-8337495, 24), to_signed(-8336067, 24), to_signed(-8334620, 24), to_signed(-8333152, 24), to_signed(-8331665, 24), to_signed(-8330159, 24), to_signed(-8328632, 24), to_signed(-8327087, 24), to_signed(-8325521, 24), to_signed(-8323936, 24), to_signed(-8322332, 24), to_signed(-8320708, 24), to_signed(-8319064, 24), to_signed(-8317401, 24), to_signed(-8315718, 24), to_signed(-8314015, 24), to_signed(-8312293, 24), to_signed(-8310552, 24), to_signed(-8308791, 24), to_signed(-8307010, 24), to_signed(-8305210, 24), to_signed(-8303390, 24), to_signed(-8301551, 24), to_signed(-8299692, 24), to_signed(-8297813, 24), to_signed(-8295916, 24), to_signed(-8293998, 24), to_signed(-8292061, 24), to_signed(-8290105, 24), to_signed(-8288129, 24), to_signed(-8286133, 24), to_signed(-8284119, 24), to_signed(-8282084, 24), to_signed(-8280030, 24), to_signed(-8277957, 24), to_signed(-8275864, 24), to_signed(-8273751, 24), to_signed(-8271620, 24), to_signed(-8269468, 24), to_signed(-8267298, 24), to_signed(-8265107, 24), to_signed(-8262898, 24), to_signed(-8260669, 24), to_signed(-8258420, 24), to_signed(-8256152, 24), to_signed(-8253865, 24), to_signed(-8251558, 24), to_signed(-8249232, 24), to_signed(-8246886, 24), to_signed(-8244521, 24), to_signed(-8242137, 24), to_signed(-8239733, 24), to_signed(-8237309, 24), to_signed(-8234867, 24), to_signed(-8232405, 24), to_signed(-8229923, 24), to_signed(-8227423, 24), to_signed(-8224903, 24), to_signed(-8222363, 24), to_signed(-8219804, 24), to_signed(-8217226, 24), to_signed(-8214629, 24), to_signed(-8212012, 24), to_signed(-8209376, 24), to_signed(-8206720, 24), to_signed(-8204046, 24), to_signed(-8201352, 24), to_signed(-8198638, 24), to_signed(-8195906, 24), to_signed(-8193154, 24), to_signed(-8190382, 24), to_signed(-8187592, 24), to_signed(-8184782, 24), to_signed(-8181953, 24), to_signed(-8179105, 24), to_signed(-8176237, 24), to_signed(-8173351, 24), to_signed(-8170445, 24), to_signed(-8167519, 24), to_signed(-8164575, 24), to_signed(-8161611, 24), to_signed(-8158629, 24), to_signed(-8155626, 24), to_signed(-8152605, 24), to_signed(-8149565, 24), to_signed(-8146505, 24), to_signed(-8143426, 24), to_signed(-8140329, 24), to_signed(-8137211, 24), to_signed(-8134075, 24), to_signed(-8130920, 24), to_signed(-8127745, 24), to_signed(-8124552, 24), to_signed(-8121339, 24), to_signed(-8118107, 24), to_signed(-8114856, 24), to_signed(-8111586, 24), to_signed(-8108297, 24), to_signed(-8104989, 24), to_signed(-8101661, 24), to_signed(-8098315, 24), to_signed(-8094950, 24), to_signed(-8091565, 24), to_signed(-8088162, 24), to_signed(-8084739, 24), to_signed(-8081298, 24), to_signed(-8077837, 24), to_signed(-8074357, 24), to_signed(-8070859, 24), to_signed(-8067341, 24), to_signed(-8063805, 24), to_signed(-8060249, 24), to_signed(-8056675, 24), to_signed(-8053081, 24), to_signed(-8049469, 24), to_signed(-8045837, 24), to_signed(-8042187, 24), to_signed(-8038518, 24), to_signed(-8034830, 24), to_signed(-8031123, 24), to_signed(-8027397, 24), to_signed(-8023652, 24), to_signed(-8019888, 24), to_signed(-8016106, 24), to_signed(-8012304, 24), to_signed(-8008484, 24), to_signed(-8004645, 24), to_signed(-8000787, 24), to_signed(-7996910, 24), to_signed(-7993015, 24), to_signed(-7989100, 24), to_signed(-7985167, 24), to_signed(-7981215, 24), to_signed(-7977244, 24), to_signed(-7973255, 24), to_signed(-7969246, 24), to_signed(-7965219, 24), to_signed(-7961173, 24), to_signed(-7957109, 24), to_signed(-7953026, 24), to_signed(-7948924, 24), to_signed(-7944803, 24), to_signed(-7940663, 24), to_signed(-7936505, 24), to_signed(-7932329, 24), to_signed(-7928133, 24), to_signed(-7923919, 24), to_signed(-7919686, 24), to_signed(-7915435, 24), to_signed(-7911165, 24), to_signed(-7906877, 24), to_signed(-7902569, 24), to_signed(-7898244, 24), to_signed(-7893899, 24), to_signed(-7889536, 24), to_signed(-7885155, 24), to_signed(-7880755, 24), to_signed(-7876336, 24), to_signed(-7871899, 24), to_signed(-7867443, 24), to_signed(-7862969, 24), to_signed(-7858476, 24), to_signed(-7853965, 24), to_signed(-7849436, 24), to_signed(-7844887, 24), to_signed(-7840321, 24), to_signed(-7835736, 24), to_signed(-7831132, 24), to_signed(-7826510, 24), to_signed(-7821870, 24), to_signed(-7817211, 24), to_signed(-7812534, 24), to_signed(-7807839, 24), to_signed(-7803125, 24), to_signed(-7798393, 24), to_signed(-7793642, 24), to_signed(-7788873, 24), to_signed(-7784086, 24), to_signed(-7779280, 24), to_signed(-7774456, 24), to_signed(-7769614, 24), to_signed(-7764754, 24), to_signed(-7759875, 24), to_signed(-7754978, 24), to_signed(-7750063, 24), to_signed(-7745129, 24), to_signed(-7740178, 24), to_signed(-7735208, 24), to_signed(-7730220, 24), to_signed(-7725213, 24), to_signed(-7720189, 24), to_signed(-7715146, 24), to_signed(-7710085, 24), to_signed(-7705006, 24), to_signed(-7699909, 24), to_signed(-7694794, 24), to_signed(-7689661, 24), to_signed(-7684509, 24), to_signed(-7679340, 24), to_signed(-7674152, 24), to_signed(-7668947, 24), to_signed(-7663723, 24), to_signed(-7658481, 24), to_signed(-7653222, 24), to_signed(-7647944, 24), to_signed(-7642648, 24), to_signed(-7637335, 24), to_signed(-7632003, 24), to_signed(-7626653, 24), to_signed(-7621286, 24), to_signed(-7615900, 24), to_signed(-7610497, 24), to_signed(-7605075, 24), to_signed(-7599636, 24), to_signed(-7594179, 24), to_signed(-7588704, 24), to_signed(-7583211, 24), to_signed(-7577701, 24), to_signed(-7572172, 24), to_signed(-7566626, 24), to_signed(-7561062, 24), to_signed(-7555480, 24), to_signed(-7549880, 24), to_signed(-7544263, 24), to_signed(-7538627, 24), to_signed(-7532974, 24), to_signed(-7527304, 24), to_signed(-7521615, 24), to_signed(-7515909, 24), to_signed(-7510185, 24), to_signed(-7504444, 24), to_signed(-7498685, 24), to_signed(-7492908, 24), to_signed(-7487114, 24), to_signed(-7481302, 24), to_signed(-7475472, 24), to_signed(-7469625, 24), to_signed(-7463760, 24), to_signed(-7457878, 24), to_signed(-7451978, 24), to_signed(-7446060, 24), to_signed(-7440125, 24), to_signed(-7434173, 24), to_signed(-7428203, 24), to_signed(-7422216, 24), to_signed(-7416211, 24), to_signed(-7410188, 24), to_signed(-7404148, 24), to_signed(-7398091, 24), to_signed(-7392017, 24), to_signed(-7385925, 24), to_signed(-7379815, 24), to_signed(-7373688, 24), to_signed(-7367544, 24), to_signed(-7361383, 24), to_signed(-7355204, 24), to_signed(-7349008, 24), to_signed(-7342795, 24), to_signed(-7336564, 24), to_signed(-7330316, 24), to_signed(-7324051, 24), to_signed(-7317769, 24), to_signed(-7311469, 24), to_signed(-7305152, 24), to_signed(-7298818, 24), to_signed(-7292467, 24), to_signed(-7286099, 24), to_signed(-7279713, 24), to_signed(-7273311, 24), to_signed(-7266891, 24), to_signed(-7260454, 24), to_signed(-7254000, 24), to_signed(-7247529, 24), to_signed(-7241041, 24), to_signed(-7234536, 24), to_signed(-7228014, 24), to_signed(-7221475, 24), to_signed(-7214919, 24), to_signed(-7208346, 24), to_signed(-7201756, 24), to_signed(-7195149, 24), to_signed(-7188525, 24), to_signed(-7181884, 24), to_signed(-7175226, 24), to_signed(-7168551, 24), to_signed(-7161860, 24), to_signed(-7155152, 24), to_signed(-7148426, 24), to_signed(-7141684, 24), to_signed(-7134926, 24), to_signed(-7128150, 24), to_signed(-7121358, 24), to_signed(-7114549, 24), to_signed(-7107723, 24), to_signed(-7100880, 24), to_signed(-7094021, 24), to_signed(-7087145, 24), to_signed(-7080252, 24), to_signed(-7073343, 24), to_signed(-7066417, 24), to_signed(-7059474, 24), to_signed(-7052515, 24), to_signed(-7045539, 24), to_signed(-7038547, 24), to_signed(-7031538, 24), to_signed(-7024512, 24), to_signed(-7017470, 24), to_signed(-7010412, 24), to_signed(-7003337, 24), to_signed(-6996245, 24), to_signed(-6989137, 24), to_signed(-6982013, 24), to_signed(-6974872, 24), to_signed(-6967715, 24), to_signed(-6960541, 24), to_signed(-6953351, 24), to_signed(-6946145, 24), to_signed(-6938922, 24), to_signed(-6931683, 24), to_signed(-6924428, 24), to_signed(-6917156, 24), to_signed(-6909868, 24), to_signed(-6902564, 24), to_signed(-6895243, 24), to_signed(-6887907, 24), to_signed(-6880554, 24), to_signed(-6873185, 24), to_signed(-6865799, 24), to_signed(-6858398, 24), to_signed(-6850980, 24), to_signed(-6843547, 24), to_signed(-6836097, 24), to_signed(-6828631, 24), to_signed(-6821149, 24), to_signed(-6813651, 24), to_signed(-6806137, 24), to_signed(-6798607, 24), to_signed(-6791061, 24), to_signed(-6783499, 24), to_signed(-6775921, 24), to_signed(-6768327, 24), to_signed(-6760718, 24), to_signed(-6753092, 24), to_signed(-6745450, 24), to_signed(-6737793, 24), to_signed(-6730119, 24), to_signed(-6722430, 24), to_signed(-6714725, 24), to_signed(-6707004, 24), to_signed(-6699268, 24), to_signed(-6691515, 24), to_signed(-6683747, 24), to_signed(-6675963, 24), to_signed(-6668164, 24), to_signed(-6660349, 24), to_signed(-6652518, 24), to_signed(-6644671, 24), to_signed(-6636809, 24), to_signed(-6628931, 24), to_signed(-6621038, 24), to_signed(-6613129, 24), to_signed(-6605204, 24), to_signed(-6597264, 24), to_signed(-6589308, 24), to_signed(-6581337, 24), to_signed(-6573351, 24), to_signed(-6565349, 24), to_signed(-6557331, 24), to_signed(-6549298, 24), to_signed(-6541250, 24), to_signed(-6533186, 24), to_signed(-6525107, 24), to_signed(-6517012, 24), to_signed(-6508902, 24), to_signed(-6500777, 24), to_signed(-6492637, 24), to_signed(-6484481, 24), to_signed(-6476310, 24), to_signed(-6468124, 24), to_signed(-6459923, 24), to_signed(-6451706, 24), to_signed(-6443474, 24), to_signed(-6435227, 24), to_signed(-6426965, 24), to_signed(-6418688, 24), to_signed(-6410395, 24), to_signed(-6402088, 24), to_signed(-6393765, 24), to_signed(-6385428, 24), to_signed(-6377075, 24), to_signed(-6368708, 24), to_signed(-6360325, 24), to_signed(-6351928, 24), to_signed(-6343515, 24), to_signed(-6335088, 24), to_signed(-6326646, 24), to_signed(-6318188, 24), to_signed(-6309716, 24), to_signed(-6301229, 24), to_signed(-6292728, 24), to_signed(-6284211, 24), to_signed(-6275680, 24), to_signed(-6267134, 24), to_signed(-6258573, 24), to_signed(-6249997, 24), to_signed(-6241407, 24), to_signed(-6232802, 24), to_signed(-6224182, 24), to_signed(-6215548, 24), to_signed(-6206899, 24), to_signed(-6198236, 24), to_signed(-6189558, 24), to_signed(-6180865, 24), to_signed(-6172158, 24), to_signed(-6163436, 24), to_signed(-6154700, 24), to_signed(-6145949, 24), to_signed(-6137184, 24), to_signed(-6128404, 24), to_signed(-6119610, 24), to_signed(-6110802, 24), to_signed(-6101979, 24), to_signed(-6093142, 24), to_signed(-6084290, 24), to_signed(-6075424, 24), to_signed(-6066544, 24), to_signed(-6057650, 24), to_signed(-6048741, 24), to_signed(-6039818, 24), to_signed(-6030881, 24), to_signed(-6021930, 24), to_signed(-6012964, 24), to_signed(-6003985, 24), to_signed(-5994991, 24), to_signed(-5985983, 24), to_signed(-5976961, 24), to_signed(-5967925, 24), to_signed(-5958875, 24), to_signed(-5949811, 24), to_signed(-5940733, 24), to_signed(-5931641, 24), to_signed(-5922535, 24), to_signed(-5913415, 24), to_signed(-5904281, 24), to_signed(-5895134, 24), to_signed(-5885972, 24), to_signed(-5876796, 24), to_signed(-5867607, 24), to_signed(-5858404, 24), to_signed(-5849187, 24), to_signed(-5839957, 24), to_signed(-5830712, 24), to_signed(-5821454, 24), to_signed(-5812182, 24), to_signed(-5802897, 24), to_signed(-5793598, 24), to_signed(-5784285, 24), to_signed(-5774958, 24), to_signed(-5765618, 24), to_signed(-5756265, 24), to_signed(-5746898, 24), to_signed(-5737517, 24), to_signed(-5728123, 24), to_signed(-5718716, 24), to_signed(-5709294, 24), to_signed(-5699860, 24), to_signed(-5690412, 24), to_signed(-5680951, 24), to_signed(-5671476, 24), to_signed(-5661988, 24), to_signed(-5652487, 24), to_signed(-5642972, 24), to_signed(-5633444, 24), to_signed(-5623903, 24), to_signed(-5614349, 24), to_signed(-5604781, 24), to_signed(-5595200, 24), to_signed(-5585606, 24), to_signed(-5575999, 24), to_signed(-5566379, 24), to_signed(-5556746, 24), to_signed(-5547099, 24), to_signed(-5537440, 24), to_signed(-5527767, 24), to_signed(-5518082, 24), to_signed(-5508384, 24), to_signed(-5498672, 24), to_signed(-5488948, 24), to_signed(-5479210, 24), to_signed(-5469460, 24), to_signed(-5459697, 24), to_signed(-5449921, 24), to_signed(-5440133, 24), to_signed(-5430331, 24), to_signed(-5420517, 24), to_signed(-5410690, 24), to_signed(-5400850, 24), to_signed(-5390997, 24), to_signed(-5381132, 24), to_signed(-5371254, 24), to_signed(-5361364, 24), to_signed(-5351461, 24), to_signed(-5341545, 24), to_signed(-5331617, 24), to_signed(-5321676, 24), to_signed(-5311723, 24), to_signed(-5301757, 24), to_signed(-5291779, 24), to_signed(-5281788, 24), to_signed(-5271785, 24), to_signed(-5261769, 24), to_signed(-5251741, 24), to_signed(-5241701, 24), to_signed(-5231648, 24), to_signed(-5221583, 24), to_signed(-5211506, 24), to_signed(-5201416, 24), to_signed(-5191315, 24), to_signed(-5181201, 24), to_signed(-5171074, 24), to_signed(-5160936, 24), to_signed(-5150786, 24), to_signed(-5140623, 24), to_signed(-5130448, 24), to_signed(-5120262, 24), to_signed(-5110063, 24), to_signed(-5099852, 24), to_signed(-5089629, 24), to_signed(-5079394, 24), to_signed(-5069147, 24), to_signed(-5058889, 24), to_signed(-5048618, 24), to_signed(-5038336, 24), to_signed(-5028041, 24), to_signed(-5017735, 24), to_signed(-5007417, 24), to_signed(-4997087, 24), to_signed(-4986746, 24), to_signed(-4976393, 24), to_signed(-4966028, 24), to_signed(-4955651, 24), to_signed(-4945263, 24), to_signed(-4934863, 24), to_signed(-4924451, 24), to_signed(-4914028, 24), to_signed(-4903593, 24), to_signed(-4893147, 24), to_signed(-4882689, 24), to_signed(-4872220, 24), to_signed(-4861739, 24), to_signed(-4851247, 24), to_signed(-4840744, 24), to_signed(-4830229, 24), to_signed(-4819702, 24), to_signed(-4809165, 24), to_signed(-4798616, 24), to_signed(-4788055, 24), to_signed(-4777484, 24), to_signed(-4766901, 24), to_signed(-4756307, 24), to_signed(-4745702, 24), to_signed(-4735086, 24), to_signed(-4724458, 24), to_signed(-4713819, 24), to_signed(-4703170, 24), to_signed(-4692509, 24), to_signed(-4681837, 24), to_signed(-4671154, 24), to_signed(-4660460, 24), to_signed(-4649756, 24), to_signed(-4639040, 24), to_signed(-4628313, 24), to_signed(-4617576, 24), to_signed(-4606827, 24), to_signed(-4596068, 24), to_signed(-4585298, 24), to_signed(-4574517, 24), to_signed(-4563725, 24), to_signed(-4552923, 24), to_signed(-4542110, 24), to_signed(-4531286, 24), to_signed(-4520452, 24), to_signed(-4509607, 24), to_signed(-4498751, 24), to_signed(-4487885, 24), to_signed(-4477008, 24), to_signed(-4466121, 24), to_signed(-4455223, 24), to_signed(-4444314, 24), to_signed(-4433396, 24), to_signed(-4422466, 24), to_signed(-4411527, 24), to_signed(-4400577, 24), to_signed(-4389616, 24), to_signed(-4378646, 24), to_signed(-4367665, 24), to_signed(-4356673, 24), to_signed(-4345672, 24), to_signed(-4334660, 24), to_signed(-4323638, 24), to_signed(-4312606, 24), to_signed(-4301564, 24), to_signed(-4290511, 24), to_signed(-4279449, 24), to_signed(-4268376, 24), to_signed(-4257293, 24), to_signed(-4246201, 24), to_signed(-4235098, 24), to_signed(-4223986, 24), to_signed(-4212863, 24), to_signed(-4201731, 24), to_signed(-4190588, 24), to_signed(-4179436, 24), to_signed(-4168274, 24), to_signed(-4157102, 24), to_signed(-4145921, 24), to_signed(-4134729, 24), to_signed(-4123528, 24), to_signed(-4112317, 24), to_signed(-4101097, 24), to_signed(-4089867, 24), to_signed(-4078627, 24), to_signed(-4067378, 24), to_signed(-4056119, 24), to_signed(-4044850, 24), to_signed(-4033572, 24), to_signed(-4022285, 24), to_signed(-4010988, 24), to_signed(-3999681, 24), to_signed(-3988366, 24), to_signed(-3977040, 24), to_signed(-3965706, 24), to_signed(-3954362, 24), to_signed(-3943009, 24), to_signed(-3931646, 24), to_signed(-3920275, 24), to_signed(-3908894, 24), to_signed(-3897504, 24), to_signed(-3886104, 24), to_signed(-3874696, 24), to_signed(-3863278, 24), to_signed(-3851852, 24), to_signed(-3840416, 24), to_signed(-3828971, 24), to_signed(-3817517, 24), to_signed(-3806055, 24), to_signed(-3794583, 24), to_signed(-3783102, 24), to_signed(-3771613, 24), to_signed(-3760114, 24), to_signed(-3748607, 24), to_signed(-3737091, 24), to_signed(-3725566, 24), to_signed(-3714032, 24), to_signed(-3702490, 24), to_signed(-3690939, 24), to_signed(-3679379, 24), to_signed(-3667811, 24), to_signed(-3656234, 24), to_signed(-3644648, 24), to_signed(-3633054, 24), to_signed(-3621451, 24), to_signed(-3609840, 24), to_signed(-3598220, 24), to_signed(-3586592, 24), to_signed(-3574955, 24), to_signed(-3563310, 24), to_signed(-3551656, 24), to_signed(-3539994, 24), to_signed(-3528324, 24), to_signed(-3516646, 24), to_signed(-3504959, 24), to_signed(-3493264, 24), to_signed(-3481561, 24), to_signed(-3469849, 24), to_signed(-3458130, 24), to_signed(-3446402, 24), to_signed(-3434666, 24), to_signed(-3422922, 24), to_signed(-3411170, 24), to_signed(-3399410, 24), to_signed(-3387642, 24), to_signed(-3375866, 24), to_signed(-3364082, 24), to_signed(-3352290, 24), to_signed(-3340491, 24), to_signed(-3328683, 24), to_signed(-3316868, 24), to_signed(-3305044, 24), to_signed(-3293213, 24), to_signed(-3281375, 24), to_signed(-3269528, 24), to_signed(-3257674, 24), to_signed(-3245812, 24), to_signed(-3233943, 24), to_signed(-3222065, 24), to_signed(-3210181, 24), to_signed(-3198289, 24), to_signed(-3186389, 24), to_signed(-3174482, 24), to_signed(-3162567, 24), to_signed(-3150645, 24), to_signed(-3138715, 24), to_signed(-3126778, 24), to_signed(-3114834, 24), to_signed(-3102882, 24), to_signed(-3090923, 24), to_signed(-3078957, 24), to_signed(-3066984, 24), to_signed(-3055003, 24), to_signed(-3043015, 24), to_signed(-3031020, 24), to_signed(-3019018, 24), to_signed(-3007009, 24), to_signed(-2994992, 24), to_signed(-2982969, 24), to_signed(-2970938, 24), to_signed(-2958901, 24), to_signed(-2946857, 24), to_signed(-2934805, 24), to_signed(-2922747, 24), to_signed(-2910682, 24), to_signed(-2898610, 24), to_signed(-2886531, 24), to_signed(-2874446, 24), to_signed(-2862354, 24), to_signed(-2850255, 24), to_signed(-2838149, 24), to_signed(-2826036, 24), to_signed(-2813917, 24), to_signed(-2801792, 24), to_signed(-2789659, 24), to_signed(-2777521, 24), to_signed(-2765375, 24), to_signed(-2753223, 24), to_signed(-2741065, 24), to_signed(-2728900, 24), to_signed(-2716729, 24), to_signed(-2704551, 24), to_signed(-2692367, 24), to_signed(-2680177, 24), to_signed(-2667980, 24), to_signed(-2655777, 24), to_signed(-2643568, 24), to_signed(-2631353, 24), to_signed(-2619131, 24), to_signed(-2606903, 24), to_signed(-2594669, 24), to_signed(-2582429, 24), to_signed(-2570183, 24), to_signed(-2557931, 24), to_signed(-2545673, 24), to_signed(-2533409, 24), to_signed(-2521139, 24), to_signed(-2508863, 24), to_signed(-2496581, 24), to_signed(-2484293, 24), to_signed(-2472000, 24), to_signed(-2459700, 24), to_signed(-2447395, 24), to_signed(-2435084, 24), to_signed(-2422767, 24), to_signed(-2410445, 24), to_signed(-2398117, 24), to_signed(-2385783, 24), to_signed(-2373443, 24), to_signed(-2361099, 24), to_signed(-2348748, 24), to_signed(-2336392, 24), to_signed(-2324030, 24), to_signed(-2311663, 24), to_signed(-2299291, 24), to_signed(-2286913, 24), to_signed(-2274530, 24), to_signed(-2262141, 24), to_signed(-2249747, 24), to_signed(-2237348, 24), to_signed(-2224944, 24), to_signed(-2212534, 24), to_signed(-2200119, 24), to_signed(-2187699, 24), to_signed(-2175274, 24), to_signed(-2162844, 24), to_signed(-2150408, 24), to_signed(-2137968, 24), to_signed(-2125522, 24), to_signed(-2113072, 24), to_signed(-2100616, 24), to_signed(-2088156, 24), to_signed(-2075690, 24), to_signed(-2063220, 24), to_signed(-2050745, 24), to_signed(-2038265, 24), to_signed(-2025780, 24), to_signed(-2013291, 24), to_signed(-2000797, 24), to_signed(-1988298, 24), to_signed(-1975794, 24), to_signed(-1963286, 24), to_signed(-1950773, 24), to_signed(-1938255, 24), to_signed(-1925733, 24), to_signed(-1913207, 24), to_signed(-1900676, 24), to_signed(-1888140, 24), to_signed(-1875600, 24), to_signed(-1863056, 24), to_signed(-1850507, 24), to_signed(-1837954, 24), to_signed(-1825396, 24), to_signed(-1812835, 24), to_signed(-1800269, 24), to_signed(-1787698, 24), to_signed(-1775124, 24), to_signed(-1762545, 24), to_signed(-1749963, 24), to_signed(-1737376, 24), to_signed(-1724785, 24), to_signed(-1712190, 24), to_signed(-1699591, 24), to_signed(-1686987, 24), to_signed(-1674380, 24), to_signed(-1661769, 24), to_signed(-1649155, 24), to_signed(-1636536, 24), to_signed(-1623913, 24), to_signed(-1611287, 24), to_signed(-1598656, 24), to_signed(-1586022, 24), to_signed(-1573385, 24), to_signed(-1560743, 24), to_signed(-1548098, 24), to_signed(-1535449, 24), to_signed(-1522797, 24), to_signed(-1510141, 24), to_signed(-1497482, 24), to_signed(-1484819, 24), to_signed(-1472152, 24), to_signed(-1459482, 24), to_signed(-1446809, 24), to_signed(-1434132, 24), to_signed(-1421452, 24), to_signed(-1408768, 24), to_signed(-1396081, 24), to_signed(-1383391, 24), to_signed(-1370698, 24), to_signed(-1358001, 24), to_signed(-1345301, 24), to_signed(-1332598, 24), to_signed(-1319892, 24), to_signed(-1307183, 24), to_signed(-1294471, 24), to_signed(-1281755, 24), to_signed(-1269037, 24), to_signed(-1256315, 24), to_signed(-1243591, 24), to_signed(-1230864, 24), to_signed(-1218134, 24), to_signed(-1205401, 24), to_signed(-1192665, 24), to_signed(-1179926, 24), to_signed(-1167185, 24), to_signed(-1154441, 24), to_signed(-1141694, 24), to_signed(-1128944, 24), to_signed(-1116192, 24), to_signed(-1103437, 24), to_signed(-1090680, 24), to_signed(-1077920, 24), to_signed(-1065157, 24), to_signed(-1052392, 24), to_signed(-1039625, 24), to_signed(-1026855, 24), to_signed(-1014082, 24), to_signed(-1001307, 24), to_signed(-988530, 24), to_signed(-975751, 24), to_signed(-962969, 24), to_signed(-950185, 24), to_signed(-937399, 24), to_signed(-924610, 24), to_signed(-911820, 24), to_signed(-899027, 24), to_signed(-886232, 24), to_signed(-873435, 24), to_signed(-860636, 24), to_signed(-847835, 24), to_signed(-835032, 24), to_signed(-822227, 24), to_signed(-809420, 24), to_signed(-796611, 24), to_signed(-783800, 24), to_signed(-770988, 24), to_signed(-758173, 24), to_signed(-745357, 24), to_signed(-732539, 24), to_signed(-719720, 24), to_signed(-706898, 24), to_signed(-694075, 24), to_signed(-681250, 24), to_signed(-668424, 24), to_signed(-655596, 24), to_signed(-642767, 24), to_signed(-629936, 24), to_signed(-617104, 24), to_signed(-604270, 24), to_signed(-591435, 24), to_signed(-578598, 24), to_signed(-565760, 24), to_signed(-552921, 24), to_signed(-540080, 24), to_signed(-527238, 24), to_signed(-514395, 24), to_signed(-501551, 24), to_signed(-488705, 24), to_signed(-475859, 24), to_signed(-463011, 24), to_signed(-450162, 24), to_signed(-437312, 24), to_signed(-424461, 24), to_signed(-411609, 24), to_signed(-398756, 24), to_signed(-385902, 24), to_signed(-373047, 24), to_signed(-360192, 24), to_signed(-347335, 24), to_signed(-334478, 24), to_signed(-321620, 24), to_signed(-308761, 24), to_signed(-295901, 24), to_signed(-283041, 24), to_signed(-270180, 24), to_signed(-257318, 24), to_signed(-244456, 24), to_signed(-231593, 24), to_signed(-218730, 24), to_signed(-205866, 24), to_signed(-193002, 24), to_signed(-180137, 24), to_signed(-167272, 24), to_signed(-154406, 24), to_signed(-141540, 24), to_signed(-128674, 24), to_signed(-115807, 24), to_signed(-102941, 24), to_signed(-90074, 24), to_signed(-77206, 24), to_signed(-64339, 24), to_signed(-51471, 24), to_signed(-38603, 24), to_signed(-25735, 24), to_signed(-12867, 24)
);
end sinewave;
