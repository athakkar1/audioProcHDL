
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library WORK;
USE work.arraypkg.ALL;

package sinewave is
  constant wave : mem := (
2047, 2068, 2090, 2111, 2133, 2154, 2175, 2197, 2218, 2239, 2261, 2282, 2303, 2324, 2346, 2367, 2388, 2409, 2430, 2451, 2472, 2493, 2514, 2535, 2555, 2576, 2597, 2617, 2638, 2658, 2679, 2699, 2719, 2739, 2759, 2779, 2799, 2819, 2839, 2858, 2878, 2897, 2917, 2936, 2955, 2974, 2993, 3012, 3031, 3050, 3068, 3087, 3105, 3123, 3141, 3159, 3177, 3195, 3212, 3230, 3247, 3264, 3281, 3298, 3315, 3331, 3348, 3364, 3380, 3396, 3412, 3428, 3444, 3459, 3474, 3489, 3504, 3519, 3534, 3548, 3563, 3577, 3591, 3604, 3618, 3632, 3645, 3658, 3671, 3684, 3696, 3709, 3721, 3733, 3745, 3756, 3768, 3779, 3790, 3801, 3812, 3823, 3833, 3843, 3853, 3863, 3872, 3882, 3891, 3900, 3909, 3917, 3926, 3934, 3942, 3950, 3957, 3965, 3972, 3979, 3986, 3992, 3999, 4005, 4011, 4017, 4022, 4028, 4033, 4038, 4042, 4047, 4051, 4055, 4059, 4063, 4067, 4070, 4073, 4076, 4078, 4081, 4083, 4085, 4087, 4089, 4090, 4091, 4092, 4093, 4094, 4094, 4094, 4095, 4094, 4094, 4093, 4093, 4092, 4090, 4089, 4087, 4086, 4084, 4081, 4079, 4076, 4074, 4071, 4067, 4064, 4061, 4057, 4053, 4049, 4045, 4040, 4035, 4031, 4026, 4020, 4015, 4009, 4004, 3998, 3992, 3985, 3979, 3972, 3966, 3959, 3952, 3944, 3937, 3929, 3921, 3913, 3905, 3897, 3889, 3880, 3872, 3863, 3854, 3844, 3835, 3826, 3816, 3806, 3797, 3787, 3776, 3766, 3756, 3745, 3735, 3724, 3713, 3702, 3691, 3679, 3668, 3656, 3645, 3633, 3621, 3609, 3597, 3585, 3573, 3560, 3548, 3535, 3523, 3510, 3497, 3484, 3471, 3458, 3445, 3432, 3418, 3405, 3391, 3378, 3364, 3350, 3337, 3323, 3309, 3295, 3281, 3267, 3253, 3239, 3225, 3210, 3196, 3182, 3167, 3153, 3138, 3124, 3109, 3095, 3080, 3066, 3051, 3036, 3022, 3007, 2992, 2978, 2963, 2948, 2934, 2919, 2904, 2889, 2875, 2860, 2845, 2831, 2816, 2801, 2787, 2772, 2757, 2743, 2728, 2714, 2699, 2685, 2670, 2656, 2641, 2627, 2613, 2598, 2584, 2570, 2556, 2542, 2528, 2514, 2500, 2486, 2472, 2459, 2445, 2431, 2418, 2404, 2391, 2378, 2364, 2351, 2338, 2325, 2312, 2299, 2286, 2274, 2261, 2249, 2236, 2224, 2212, 2199, 2187, 2175, 2163, 2152, 2140, 2128, 2117, 2106, 2094, 2083, 2072, 2061, 2051, 2040, 2029, 2019, 2009, 1998, 1988, 1978, 1968, 1959, 1949, 1940, 1930, 1921, 1912, 1903, 1894, 1885, 1877, 1868, 1860, 1852, 1844, 1836, 1828, 1820, 1813, 1805, 1798, 1791, 1784, 1777, 1770, 1764, 1758, 1751, 1745, 1739, 1733, 1728, 1722, 1717, 1711, 1706, 1701, 1696, 1692, 1687, 1683, 1679, 1675, 1671, 1667, 1663, 1660, 1656, 1653, 1650, 1647, 1644, 1641, 1639, 1637, 1634, 1632, 1630, 1628, 1627, 1625, 1624, 1623, 1622, 1621, 1620, 1619, 1619, 1618, 1618, 1618, 1618, 1618, 1618, 1619, 1619, 1620, 1621, 1622, 1623, 1624, 1625, 1627, 1628, 1630, 1632, 1634, 1636, 1638, 1640, 1643, 1645, 1648, 1651, 1653, 1656, 1660, 1663, 1666, 1670, 1673, 1677, 1681, 1684, 1688, 1692, 1697, 1701, 1705, 1710, 1714, 1719, 1724, 1728, 1733, 1738, 1743, 1749, 1754, 1759, 1765, 1770, 1776, 1781, 1787, 1793, 1799, 1805, 1810, 1817, 1823, 1829, 1835, 1841, 1848, 1854, 1860, 1867, 1873, 1880, 1887, 1893, 1900, 1907, 1914, 1920, 1927, 1934, 1941, 1948, 1955, 1962, 1969, 1976, 1983, 1990, 1997, 2004, 2011, 2018, 2026, 2033, 2040, 2047, 2054, 2061, 2068, 2076, 2083, 2090, 2097, 2104, 2111, 2118, 2125, 2132, 2139, 2146, 2153, 2160, 2167, 2174, 2180, 2187, 2194, 2201, 2207, 2214, 2221, 2227, 2234, 2240, 2246, 2253, 2259, 2265, 2271, 2277, 2284, 2289, 2295, 2301, 2307, 2313, 2318, 2324, 2329, 2335, 2340, 2345, 2351, 2356, 2361, 2366, 2370, 2375, 2380, 2384, 2389, 2393, 2397, 2402, 2406, 2410, 2413, 2417, 2421, 2424, 2428, 2431, 2434, 2438, 2441, 2443, 2446, 2449, 2451, 2454, 2456, 2458, 2460, 2462, 2464, 2466, 2467, 2469, 2470, 2471, 2472, 2473, 2474, 2475, 2475, 2476, 2476, 2476, 2476, 2476, 2476, 2475, 2475, 2474, 2473, 2472, 2471, 2470, 2469, 2467, 2466, 2464, 2462, 2460, 2457, 2455, 2453, 2450, 2447, 2444, 2441, 2438, 2434, 2431, 2427, 2423, 2419, 2415, 2411, 2407, 2402, 2398, 2393, 2388, 2383, 2377, 2372, 2366, 2361, 2355, 2349, 2343, 2336, 2330, 2324, 2317, 2310, 2303, 2296, 2289, 2281, 2274, 2266, 2258, 2250, 2242, 2234, 2226, 2217, 2209, 2200, 2191, 2182, 2173, 2164, 2154, 2145, 2135, 2126, 2116, 2106, 2096, 2085, 2075, 2065, 2054, 2043, 2033, 2022, 2011, 2000, 1988, 1977, 1966, 1954, 1942, 1931, 1919, 1907, 1895, 1882, 1870, 1858, 1845, 1833, 1820, 1808, 1795, 1782, 1769, 1756, 1743, 1730, 1716, 1703, 1690, 1676, 1663, 1649, 1635, 1622, 1608, 1594, 1580, 1566, 1552, 1538, 1524, 1510, 1496, 1481, 1467, 1453, 1438, 1424, 1409, 1395, 1380, 1366, 1351, 1337, 1322, 1307, 1293, 1278, 1263, 1249, 1234, 1219, 1205, 1190, 1175, 1160, 1146, 1131, 1116, 1102, 1087, 1072, 1058, 1043, 1028, 1014, 999, 985, 970, 956, 941, 927, 912, 898, 884, 869, 855, 841, 827, 813, 799, 785, 771, 757, 744, 730, 716, 703, 689, 676, 662, 649, 636, 623, 610, 597, 584, 571, 559, 546, 534, 521, 509, 497, 485, 473, 461, 449, 438, 426, 415, 403, 392, 381, 370, 359, 349, 338, 328, 318, 307, 297, 288, 278, 268, 259, 250, 240, 231, 222, 214, 205, 197, 189, 181, 173, 165, 157, 150, 142, 135, 128, 122, 115, 109, 102, 96, 90, 85, 79, 74, 68, 63, 59, 54, 49, 45, 41, 37, 33, 30, 27, 23, 20, 18, 15, 13, 10, 8, 7, 5, 4, 2, 1, 1, 0, 0, 0, 0, 0, 0, 1, 2, 3, 4, 5, 7, 9, 11, 13, 16, 18, 21, 24, 27, 31, 35, 39, 43, 47, 52, 56, 61, 66, 72, 77, 83, 89, 95, 102, 108, 115, 122, 129, 137, 144, 152, 160, 168, 177, 185, 194, 203, 212, 222, 231, 241, 251, 261, 271, 282, 293, 304, 315, 326, 338, 349, 361, 373, 385, 398, 410, 423, 436, 449, 462, 476, 490, 503, 517, 531, 546, 560, 575, 590, 605, 620, 635, 650, 666, 682, 698, 714, 730, 746, 763, 779, 796, 813, 830, 847, 864, 882, 899, 917, 935, 953, 971, 989, 1007, 1026, 1044, 1063, 1082, 1101, 1120, 1139, 1158, 1177, 1197, 1216, 1236, 1255, 1275, 1295, 1315, 1335, 1355, 1375, 1395, 1415, 1436, 1456, 1477, 1497, 1518, 1539, 1559, 1580, 1601, 1622, 1643, 1664, 1685, 1706, 1727, 1748, 1770, 1791, 1812, 1833, 1855, 1876, 1897, 1919, 1940, 1961, 1983, 2004, 2026
);
end sinewave;
