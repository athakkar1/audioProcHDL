
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.fixed_pkg.ALL;
LIBRARY work;
USE work.arraypkg.all;
package mask_gen is
    CONSTANT decimal_numbers: mask := (
0 => to_sfixed(0.000000000000000000, mask_point'left, mask_point'right),
1 => to_sfixed(0.000000483772800220, mask_point'left, mask_point'right),
2 => to_sfixed(0.000002549496307422, mask_point'left, mask_point'right),
3 => to_sfixed(0.000004493049991311, mask_point'left, mask_point'right),
4 => to_sfixed(0.000001977300870945, mask_point'left, mask_point'right),
5 => to_sfixed(-0.000008096026285026, mask_point'left, mask_point'right),
6 => to_sfixed(-0.000022962880906526, mask_point'left, mask_point'right),
7 => to_sfixed(-0.000032668316664624, mask_point'left, mask_point'right),
8 => to_sfixed(-0.000024593942330213, mask_point'left, mask_point'right),
9 => to_sfixed(0.000007457137450783, mask_point'left, mask_point'right),
10 => to_sfixed(0.000054903489217594, mask_point'left, mask_point'right),
11 => to_sfixed(0.000093354585877513, mask_point'left, mask_point'right),
12 => to_sfixed(0.000092526144235900, mask_point'left, mask_point'right),
13 => to_sfixed(0.000034325439060294, mask_point'left, mask_point'right),
14 => to_sfixed(-0.000070145615172208, mask_point'left, mask_point'right),
15 => to_sfixed(-0.000176250008270958, mask_point'left, mask_point'right),
16 => to_sfixed(-0.000221249559833396, mask_point'left, mask_point'right),
17 => to_sfixed(-0.000156322383172309, mask_point'left, mask_point'right),
18 => to_sfixed(0.000019319209665833, mask_point'left, mask_point'right),
19 => to_sfixed(0.000242284558165956, mask_point'left, mask_point'right),
20 => to_sfixed(0.000401878818695863, mask_point'left, mask_point'right),
21 => to_sfixed(0.000389627128031404, mask_point'left, mask_point'right),
22 => to_sfixed(0.000161769974507884, mask_point'left, mask_point'right),
23 => to_sfixed(-0.000217777884892742, mask_point'left, mask_point'right),
24 => to_sfixed(-0.000583763323780547, mask_point'left, mask_point'right),
25 => to_sfixed(-0.000734436629725747, mask_point'left, mask_point'right),
26 => to_sfixed(-0.000533278213991954, mask_point'left, mask_point'right),
27 => to_sfixed(0.000000000000000005, mask_point'left, mask_point'right),
28 => to_sfixed(0.000662130951727776, mask_point'left, mask_point'right),
29 => to_sfixed(0.001132622797279600, mask_point'left, mask_point'right),
30 => to_sfixed(0.001118957008569579, mask_point'left, mask_point'right),
31 => to_sfixed(0.000519398350991118, mask_point'left, mask_point'right),
32 => to_sfixed(-0.000480760449723781, mask_point'left, mask_point'right),
33 => to_sfixed(-0.001445573839536363, mask_point'left, mask_point'right),
34 => to_sfixed(-0.001865789851114064, mask_point'left, mask_point'right),
35 => to_sfixed(-0.001411591106940711, mask_point'left, mask_point'right),
36 => to_sfixed(-0.000141735699087744, mask_point'left, mask_point'right),
37 => to_sfixed(0.001450101489474747, mask_point'left, mask_point'right),
38 => to_sfixed(0.002607743145481599, mask_point'left, mask_point'right),
39 => to_sfixed(0.002654807280008334, mask_point'left, mask_point'right),
40 => to_sfixed(0.001359627210756587, mask_point'left, mask_point'right),
41 => to_sfixed(-0.000863229674027558, mask_point'left, mask_point'right),
42 => to_sfixed(-0.003049021318228376, mask_point'left, mask_point'right),
43 => to_sfixed(-0.004079604946561900, mask_point'left, mask_point'right),
44 => to_sfixed(-0.003228746056077710, mask_point'left, mask_point'right),
45 => to_sfixed(-0.000600972698884819, mask_point'left, mask_point'right),
46 => to_sfixed(0.002779267078060167, mask_point'left, mask_point'right),
47 => to_sfixed(0.005332423361351708, mask_point'left, mask_point'right),
48 => to_sfixed(0.005631804466623587, mask_point'left, mask_point'right),
49 => to_sfixed(0.003150856937418233, mask_point'left, mask_point'right),
50 => to_sfixed(-0.001322809024486645, mask_point'left, mask_point'right),
51 => to_sfixed(-0.005869525897873455, mask_point'left, mask_point'right),
52 => to_sfixed(-0.008218950341616701, mask_point'left, mask_point'right),
53 => to_sfixed(-0.006832710381255036, mask_point'left, mask_point'right),
54 => to_sfixed(-0.001793109131179641, mask_point'left, mask_point'right),
55 => to_sfixed(0.004976445608570192, mask_point'left, mask_point'right),
56 => to_sfixed(0.010373300679926933, mask_point'left, mask_point'right),
57 => to_sfixed(0.011468700024768028, mask_point'left, mask_point'right),
58 => to_sfixed(0.006990930317331622, mask_point'left, mask_point'right),
59 => to_sfixed(-0.001771481509888936, mask_point'left, mask_point'right),
60 => to_sfixed(-0.011179951451509969, mask_point'left, mask_point'right),
61 => to_sfixed(-0.016641911929546845, mask_point'left, mask_point'right),
62 => to_sfixed(-0.014703391121280518, mask_point'left, mask_point'right),
63 => to_sfixed(-0.004941117294168649, mask_point'left, mask_point'right),
64 => to_sfixed(0.009282361850304557, mask_point'left, mask_point'right),
65 => to_sfixed(0.021742338718174912, mask_point'left, mask_point'right),
66 => to_sfixed(0.025796269275013488, mask_point'left, mask_point'right),
67 => to_sfixed(0.017470754442428061, mask_point'left, mask_point'right),
68 => to_sfixed(-0.002100958650438089, mask_point'left, mask_point'right),
69 => to_sfixed(-0.026070400720082380, mask_point'left, mask_point'right),
70 => to_sfixed(-0.043627924524548188, mask_point'left, mask_point'right),
71 => to_sfixed(-0.043704593010747257, mask_point'left, mask_point'right),
72 => to_sfixed(-0.019339622962815228, mask_point'left, mask_point'right),
73 => to_sfixed(0.028976270321158695, mask_point'left, mask_point'right),
74 => to_sfixed(0.092410108993059376, mask_point'left, mask_point'right),
75 => to_sfixed(0.155910702475902579, mask_point'left, mask_point'right),
76 => to_sfixed(0.202761369724884566, mask_point'left, mask_point'right),
77 => to_sfixed(0.220001571525003131, mask_point'left, mask_point'right),
78 => to_sfixed(0.202761369724884566, mask_point'left, mask_point'right),
79 => to_sfixed(0.155910702475902579, mask_point'left, mask_point'right),
80 => to_sfixed(0.092410108993059376, mask_point'left, mask_point'right),
81 => to_sfixed(0.028976270321158695, mask_point'left, mask_point'right),
82 => to_sfixed(-0.019339622962815235, mask_point'left, mask_point'right),
83 => to_sfixed(-0.043704593010747257, mask_point'left, mask_point'right),
84 => to_sfixed(-0.043627924524548188, mask_point'left, mask_point'right),
85 => to_sfixed(-0.026070400720082380, mask_point'left, mask_point'right),
86 => to_sfixed(-0.002100958650438090, mask_point'left, mask_point'right),
87 => to_sfixed(0.017470754442428068, mask_point'left, mask_point'right),
88 => to_sfixed(0.025796269275013495, mask_point'left, mask_point'right),
89 => to_sfixed(0.021742338718174915, mask_point'left, mask_point'right),
90 => to_sfixed(0.009282361850304557, mask_point'left, mask_point'right),
91 => to_sfixed(-0.004941117294168649, mask_point'left, mask_point'right),
92 => to_sfixed(-0.014703391121280524, mask_point'left, mask_point'right),
93 => to_sfixed(-0.016641911929546848, mask_point'left, mask_point'right),
94 => to_sfixed(-0.011179951451509969, mask_point'left, mask_point'right),
95 => to_sfixed(-0.001771481509888936, mask_point'left, mask_point'right),
96 => to_sfixed(0.006990930317331622, mask_point'left, mask_point'right),
97 => to_sfixed(0.011468700024768031, mask_point'left, mask_point'right),
98 => to_sfixed(0.010373300679926938, mask_point'left, mask_point'right),
99 => to_sfixed(0.004976445608570193, mask_point'left, mask_point'right),
100 => to_sfixed(-0.001793109131179640, mask_point'left, mask_point'right),
101 => to_sfixed(-0.006832710381255036, mask_point'left, mask_point'right),
102 => to_sfixed(-0.008218950341616701, mask_point'left, mask_point'right),
103 => to_sfixed(-0.005869525897873455, mask_point'left, mask_point'right),
104 => to_sfixed(-0.001322809024486645, mask_point'left, mask_point'right),
105 => to_sfixed(0.003150856937418233, mask_point'left, mask_point'right),
106 => to_sfixed(0.005631804466623589, mask_point'left, mask_point'right),
107 => to_sfixed(0.005332423361351707, mask_point'left, mask_point'right),
108 => to_sfixed(0.002779267078060168, mask_point'left, mask_point'right),
109 => to_sfixed(-0.000600972698884819, mask_point'left, mask_point'right),
110 => to_sfixed(-0.003228746056077713, mask_point'left, mask_point'right),
111 => to_sfixed(-0.004079604946561899, mask_point'left, mask_point'right),
112 => to_sfixed(-0.003049021318228376, mask_point'left, mask_point'right),
113 => to_sfixed(-0.000863229674027559, mask_point'left, mask_point'right),
114 => to_sfixed(0.001359627210756587, mask_point'left, mask_point'right),
115 => to_sfixed(0.002654807280008333, mask_point'left, mask_point'right),
116 => to_sfixed(0.002607743145481599, mask_point'left, mask_point'right),
117 => to_sfixed(0.001450101489474749, mask_point'left, mask_point'right),
118 => to_sfixed(-0.000141735699087744, mask_point'left, mask_point'right),
119 => to_sfixed(-0.001411591106940712, mask_point'left, mask_point'right),
120 => to_sfixed(-0.001865789851114066, mask_point'left, mask_point'right),
121 => to_sfixed(-0.001445573839536364, mask_point'left, mask_point'right),
122 => to_sfixed(-0.000480760449723781, mask_point'left, mask_point'right),
123 => to_sfixed(0.000519398350991118, mask_point'left, mask_point'right),
124 => to_sfixed(0.001118957008569580, mask_point'left, mask_point'right),
125 => to_sfixed(0.001132622797279602, mask_point'left, mask_point'right),
126 => to_sfixed(0.000662130951727775, mask_point'left, mask_point'right),
127 => to_sfixed(0.000000000000000005, mask_point'left, mask_point'right),
128 => to_sfixed(-0.000533278213991955, mask_point'left, mask_point'right),
129 => to_sfixed(-0.000734436629725749, mask_point'left, mask_point'right),
130 => to_sfixed(-0.000583763323780548, mask_point'left, mask_point'right),
131 => to_sfixed(-0.000217777884892742, mask_point'left, mask_point'right),
132 => to_sfixed(0.000161769974507884, mask_point'left, mask_point'right),
133 => to_sfixed(0.000389627128031403, mask_point'left, mask_point'right),
134 => to_sfixed(0.000401878818695863, mask_point'left, mask_point'right),
135 => to_sfixed(0.000242284558165956, mask_point'left, mask_point'right),
136 => to_sfixed(0.000019319209665833, mask_point'left, mask_point'right),
137 => to_sfixed(-0.000156322383172309, mask_point'left, mask_point'right),
138 => to_sfixed(-0.000221249559833396, mask_point'left, mask_point'right),
139 => to_sfixed(-0.000176250008270959, mask_point'left, mask_point'right),
140 => to_sfixed(-0.000070145615172208, mask_point'left, mask_point'right),
141 => to_sfixed(0.000034325439060294, mask_point'left, mask_point'right),
142 => to_sfixed(0.000092526144235900, mask_point'left, mask_point'right),
143 => to_sfixed(0.000093354585877513, mask_point'left, mask_point'right),
144 => to_sfixed(0.000054903489217595, mask_point'left, mask_point'right),
145 => to_sfixed(0.000007457137450783, mask_point'left, mask_point'right),
146 => to_sfixed(-0.000024593942330213, mask_point'left, mask_point'right),
147 => to_sfixed(-0.000032668316664624, mask_point'left, mask_point'right),
148 => to_sfixed(-0.000022962880906526, mask_point'left, mask_point'right),
149 => to_sfixed(-0.000008096026285026, mask_point'left, mask_point'right),
150 => to_sfixed(0.000001977300870945, mask_point'left, mask_point'right),
151 => to_sfixed(0.000004493049991311, mask_point'left, mask_point'right),
152 => to_sfixed(0.000002549496307422, mask_point'left, mask_point'right),
153 => to_sfixed(0.000000483772800221, mask_point'left, mask_point'right),
154 => to_sfixed(0.000000000000000000, mask_point'left, mask_point'right)

);
END mask_gen;
