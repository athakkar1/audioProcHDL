
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.fixed_pkg.ALL;
LIBRARY work;
USE work.arraypkg.all;
package mask_gen is
    CONSTANT decimal_numbers: mask := (
0 => to_sfixed(0.000000000000000000, mask_point'left, mask_point'right),
1 => to_sfixed(0.000007089254541241, mask_point'left, mask_point'right),
2 => to_sfixed(0.000040982153450201, mask_point'left, mask_point'right),
3 => to_sfixed(0.000114844201775314, mask_point'left, mask_point'right),
4 => to_sfixed(0.000229282466569670, mask_point'left, mask_point'right),
5 => to_sfixed(0.000366449499768783, mask_point'left, mask_point'right),
6 => to_sfixed(0.000485554151555692, mask_point'left, mask_point'right),
7 => to_sfixed(0.000521739991755640, mask_point'left, mask_point'right),
8 => to_sfixed(0.000390575038207813, mask_point'left, mask_point'right),
9 => to_sfixed(0.000000000000000000, mask_point'left, mask_point'right),
10 => to_sfixed(-0.000729631515130406, mask_point'left, mask_point'right),
11 => to_sfixed(-0.001838720477456150, mask_point'left, mask_point'right),
12 => to_sfixed(-0.003298397915155672, mask_point'left, mask_point'right),
13 => to_sfixed(-0.004983026030425332, mask_point'left, mask_point'right),
14 => to_sfixed(-0.006652247065974609, mask_point'left, mask_point'right),
15 => to_sfixed(-0.007949546407311679, mask_point'left, mask_point'right),
16 => to_sfixed(-0.008422577180419980, mask_point'left, mask_point'right),
17 => to_sfixed(-0.007567170301013336, mask_point'left, mask_point'right),
18 => to_sfixed(-0.004892489896200722, mask_point'left, mask_point'right),
19 => to_sfixed(0.000000000000000002, mask_point'left, mask_point'right),
20 => to_sfixed(0.007335206643526098, mask_point'left, mask_point'right),
21 => to_sfixed(0.017094609576550658, mask_point'left, mask_point'right),
22 => to_sfixed(0.028971907681722187, mask_point'left, mask_point'right),
23 => to_sfixed(0.042365331159356215, mask_point'left, mask_point'right),
24 => to_sfixed(0.056412667295446355, mask_point'left, mask_point'right),
25 => to_sfixed(0.070068200301094521, mask_point'left, mask_point'right),
26 => to_sfixed(0.082213446391851713, mask_point'left, mask_point'right),
27 => to_sfixed(0.091787166614097526, mask_point'left, mask_point'right),
28 => to_sfixed(0.097915951452103259, mask_point'left, mask_point'right),
29 => to_sfixed(0.100025605831429137, mask_point'left, mask_point'right),
30 => to_sfixed(0.097915951452103259, mask_point'left, mask_point'right),
31 => to_sfixed(0.091787166614097526, mask_point'left, mask_point'right),
32 => to_sfixed(0.082213446391851713, mask_point'left, mask_point'right),
33 => to_sfixed(0.070068200301094508, mask_point'left, mask_point'right),
34 => to_sfixed(0.056412667295446355, mask_point'left, mask_point'right),
35 => to_sfixed(0.042365331159356229, mask_point'left, mask_point'right),
36 => to_sfixed(0.028971907681722201, mask_point'left, mask_point'right),
37 => to_sfixed(0.017094609576550655, mask_point'left, mask_point'right),
38 => to_sfixed(0.007335206643526100, mask_point'left, mask_point'right),
39 => to_sfixed(0.000000000000000002, mask_point'left, mask_point'right),
40 => to_sfixed(-0.004892489896200725, mask_point'left, mask_point'right),
41 => to_sfixed(-0.007567170301013340, mask_point'left, mask_point'right),
42 => to_sfixed(-0.008422577180419980, mask_point'left, mask_point'right),
43 => to_sfixed(-0.007949546407311688, mask_point'left, mask_point'right),
44 => to_sfixed(-0.006652247065974618, mask_point'left, mask_point'right),
45 => to_sfixed(-0.004983026030425335, mask_point'left, mask_point'right),
46 => to_sfixed(-0.003298397915155677, mask_point'left, mask_point'right),
47 => to_sfixed(-0.001838720477456152, mask_point'left, mask_point'right),
48 => to_sfixed(-0.000729631515130406, mask_point'left, mask_point'right),
49 => to_sfixed(0.000000000000000000, mask_point'left, mask_point'right),
50 => to_sfixed(0.000390575038207813, mask_point'left, mask_point'right),
51 => to_sfixed(0.000521739991755639, mask_point'left, mask_point'right),
52 => to_sfixed(0.000485554151555692, mask_point'left, mask_point'right),
53 => to_sfixed(0.000366449499768783, mask_point'left, mask_point'right),
54 => to_sfixed(0.000229282466569670, mask_point'left, mask_point'right),
55 => to_sfixed(0.000114844201775314, mask_point'left, mask_point'right),
56 => to_sfixed(0.000040982153450201, mask_point'left, mask_point'right),
57 => to_sfixed(0.000007089254541241, mask_point'left, mask_point'right),
58 => to_sfixed(0.000000000000000000, mask_point'left, mask_point'right)

);
END mask_gen;
