
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;
library WORK;
USE work.arraypkg.ALL;

package sinewave is
  constant wave : mem := (
to_signed(0, 24), to_signed(7967, 24), to_signed(15935, 24), to_signed(23903, 24), to_signed(31871, 24), to_signed(39839, 24), to_signed(47807, 24), to_signed(55774, 24), to_signed(63742, 24), to_signed(71709, 24), to_signed(79676, 24), to_signed(87643, 24), to_signed(95610, 24), to_signed(103576, 24), to_signed(111542, 24), to_signed(119508, 24), to_signed(127474, 24), to_signed(135440, 24), to_signed(143405, 24), to_signed(151369, 24), to_signed(159334, 24), to_signed(167298, 24), to_signed(175261, 24), to_signed(183225, 24), to_signed(191187, 24), to_signed(199150, 24), to_signed(207112, 24), to_signed(215073, 24), to_signed(223034, 24), to_signed(230994, 24), to_signed(238954, 24), to_signed(246913, 24), to_signed(254872, 24), to_signed(262830, 24), to_signed(270787, 24), to_signed(278744, 24), to_signed(286700, 24), to_signed(294656, 24), to_signed(302611, 24), to_signed(310565, 24), to_signed(318518, 24), to_signed(326471, 24), to_signed(334422, 24), to_signed(342373, 24), to_signed(350324, 24), to_signed(358273, 24), to_signed(366222, 24), to_signed(374169, 24), to_signed(382116, 24), to_signed(390062, 24), to_signed(398007, 24), to_signed(405951, 24), to_signed(413894, 24), to_signed(421836, 24), to_signed(429778, 24), to_signed(437718, 24), to_signed(445657, 24), to_signed(453595, 24), to_signed(461532, 24), to_signed(469468, 24), to_signed(477403, 24), to_signed(485336, 24), to_signed(493269, 24), to_signed(501200, 24), to_signed(509130, 24), to_signed(517059, 24), to_signed(524987, 24), to_signed(532914, 24), to_signed(540839, 24), to_signed(548763, 24), to_signed(556686, 24), to_signed(564607, 24), to_signed(572527, 24), to_signed(580446, 24), to_signed(588363, 24), to_signed(596279, 24), to_signed(604194, 24), to_signed(612107, 24), to_signed(620019, 24), to_signed(627929, 24), to_signed(635838, 24), to_signed(643745, 24), to_signed(651651, 24), to_signed(659555, 24), to_signed(667458, 24), to_signed(675359, 24), to_signed(683258, 24), to_signed(691156, 24), to_signed(699053, 24), to_signed(706947, 24), to_signed(714840, 24), to_signed(722732, 24), to_signed(730621, 24), to_signed(738509, 24), to_signed(746395, 24), to_signed(754280, 24), to_signed(762162, 24), to_signed(770043, 24), to_signed(777922, 24), to_signed(785799, 24), to_signed(793675, 24), to_signed(801548, 24), to_signed(809420, 24), to_signed(817289, 24), to_signed(825157, 24), to_signed(833023, 24), to_signed(840887, 24), to_signed(848749, 24), to_signed(856608, 24), to_signed(864466, 24), to_signed(872322, 24), to_signed(880176, 24), to_signed(888028, 24), to_signed(895877, 24), to_signed(903725, 24), to_signed(911570, 24), to_signed(919413, 24), to_signed(927254, 24), to_signed(935093, 24), to_signed(942930, 24), to_signed(950764, 24), to_signed(958597, 24), to_signed(966427, 24), to_signed(974254, 24), to_signed(982080, 24), to_signed(989903, 24), to_signed(997723, 24), to_signed(1005542, 24), to_signed(1013358, 24), to_signed(1021172, 24), to_signed(1028983, 24), to_signed(1036792, 24), to_signed(1044598, 24), to_signed(1052402, 24), to_signed(1060204, 24), to_signed(1068002, 24), to_signed(1075799, 24), to_signed(1083593, 24), to_signed(1091384, 24), to_signed(1099173, 24), to_signed(1106959, 24), to_signed(1114743, 24), to_signed(1122524, 24), to_signed(1130302, 24), to_signed(1138078, 24), to_signed(1145851, 24), to_signed(1153621, 24), to_signed(1161389, 24), to_signed(1169154, 24), to_signed(1176916, 24), to_signed(1184675, 24), to_signed(1192432, 24), to_signed(1200186, 24), to_signed(1207936, 24), to_signed(1215685, 24), to_signed(1223430, 24), to_signed(1231172, 24), to_signed(1238912, 24), to_signed(1246648, 24), to_signed(1254382, 24), to_signed(1262112, 24), to_signed(1269840, 24), to_signed(1277565, 24), to_signed(1285286, 24), to_signed(1293005, 24), to_signed(1300721, 24), to_signed(1308433, 24), to_signed(1316143, 24), to_signed(1323849, 24), to_signed(1331552, 24), to_signed(1339253, 24), to_signed(1346950, 24), to_signed(1354643, 24), to_signed(1362334, 24), to_signed(1370021, 24), to_signed(1377706, 24), to_signed(1385387, 24), to_signed(1393064, 24), to_signed(1400739, 24), to_signed(1408410, 24), to_signed(1416078, 24), to_signed(1423742, 24), to_signed(1431403, 24), to_signed(1439061, 24), to_signed(1446715, 24), to_signed(1454366, 24), to_signed(1462014, 24), to_signed(1469658, 24), to_signed(1477299, 24), to_signed(1484936, 24), to_signed(1492570, 24), to_signed(1500200, 24), to_signed(1507826, 24), to_signed(1515449, 24), to_signed(1523069, 24), to_signed(1530685, 24), to_signed(1538297, 24), to_signed(1545906, 24), to_signed(1553511, 24), to_signed(1561112, 24), to_signed(1568710, 24), to_signed(1576304, 24), to_signed(1583895, 24), to_signed(1591481, 24), to_signed(1599064, 24), to_signed(1606643, 24), to_signed(1614219, 24), to_signed(1621790, 24), to_signed(1629358, 24), to_signed(1636922, 24), to_signed(1644482, 24), to_signed(1652038, 24), to_signed(1659590, 24), to_signed(1667139, 24), to_signed(1674683, 24), to_signed(1682224, 24), to_signed(1689760, 24), to_signed(1697293, 24), to_signed(1704821, 24), to_signed(1712346, 24), to_signed(1719866, 24), to_signed(1727383, 24), to_signed(1734895, 24), to_signed(1742404, 24), to_signed(1749908, 24), to_signed(1757408, 24), to_signed(1764904, 24), to_signed(1772396, 24), to_signed(1779883, 24), to_signed(1787367, 24), to_signed(1794846, 24), to_signed(1802321, 24), to_signed(1809792, 24), to_signed(1817259, 24), to_signed(1824721, 24), to_signed(1832179, 24), to_signed(1839633, 24), to_signed(1847082, 24), to_signed(1854527, 24), to_signed(1861967, 24), to_signed(1869404, 24), to_signed(1876836, 24), to_signed(1884263, 24), to_signed(1891686, 24), to_signed(1899105, 24), to_signed(1906519, 24), to_signed(1913928, 24), to_signed(1921333, 24), to_signed(1928734, 24), to_signed(1936130, 24), to_signed(1943521, 24), to_signed(1950908, 24), to_signed(1958291, 24), to_signed(1965668, 24), to_signed(1973041, 24), to_signed(1980410, 24), to_signed(1987774, 24), to_signed(1995133, 24), to_signed(2002487, 24), to_signed(2009837, 24), to_signed(2017182, 24), to_signed(2024522, 24), to_signed(2031857, 24), to_signed(2039188, 24), to_signed(2046514, 24), to_signed(2053835, 24), to_signed(2061151, 24), to_signed(2068463, 24), to_signed(2075769, 24), to_signed(2083071, 24), to_signed(2090367, 24), to_signed(2097659, 24), to_signed(2104946, 24), to_signed(2112228, 24), to_signed(2119505, 24), to_signed(2126777, 24), to_signed(2134044, 24), to_signed(2141306, 24), to_signed(2148563, 24), to_signed(2155814, 24), to_signed(2163061, 24), to_signed(2170303, 24), to_signed(2177539, 24), to_signed(2184771, 24), to_signed(2191997, 24), to_signed(2199218, 24), to_signed(2206434, 24), to_signed(2213645, 24), to_signed(2220851, 24), to_signed(2228051, 24), to_signed(2235246, 24), to_signed(2242436, 24), to_signed(2249620, 24), to_signed(2256800, 24), to_signed(2263974, 24), to_signed(2271142, 24), to_signed(2278306, 24), to_signed(2285464, 24), to_signed(2292616, 24), to_signed(2299763, 24), to_signed(2306905, 24), to_signed(2314041, 24), to_signed(2321172, 24), to_signed(2328298, 24), to_signed(2335417, 24), to_signed(2342532, 24), to_signed(2349641, 24), to_signed(2356744, 24), to_signed(2363842, 24), to_signed(2370934, 24), to_signed(2378021, 24), to_signed(2385102, 24), to_signed(2392178, 24), to_signed(2399247, 24), to_signed(2406312, 24), to_signed(2413370, 24), to_signed(2420423, 24), to_signed(2427470, 24), to_signed(2434512, 24), to_signed(2441547, 24), to_signed(2448577, 24), to_signed(2455602, 24), to_signed(2462620, 24), to_signed(2469633, 24), to_signed(2476640, 24), to_signed(2483641, 24), to_signed(2490636, 24), to_signed(2497625, 24), to_signed(2504609, 24), to_signed(2511586, 24), to_signed(2518558, 24), to_signed(2525523, 24), to_signed(2532483, 24), to_signed(2539437, 24), to_signed(2546385, 24), to_signed(2553327, 24), to_signed(2560263, 24), to_signed(2567192, 24), to_signed(2574116, 24), to_signed(2581034, 24), to_signed(2587945, 24), to_signed(2594851, 24), to_signed(2601750, 24), to_signed(2608644, 24), to_signed(2615531, 24), to_signed(2622412, 24), to_signed(2629287, 24), to_signed(2636155, 24), to_signed(2643018, 24), to_signed(2649874, 24), to_signed(2656724, 24), to_signed(2663568, 24), to_signed(2670405, 24), to_signed(2677237, 24), to_signed(2684062, 24), to_signed(2690880, 24), to_signed(2697692, 24), to_signed(2704498, 24), to_signed(2711298, 24), to_signed(2718091, 24), to_signed(2724878, 24), to_signed(2731658, 24), to_signed(2738432, 24), to_signed(2745200, 24), to_signed(2751961, 24), to_signed(2758715, 24), to_signed(2765463, 24), to_signed(2772205, 24), to_signed(2778940, 24), to_signed(2785668, 24), to_signed(2792390, 24), to_signed(2799106, 24), to_signed(2805814, 24), to_signed(2812517, 24), to_signed(2819212, 24), to_signed(2825901, 24), to_signed(2832583, 24), to_signed(2839259, 24), to_signed(2845928, 24), to_signed(2852590, 24), to_signed(2859246, 24), to_signed(2865894, 24), to_signed(2872536, 24), to_signed(2879172, 24), to_signed(2885800, 24), to_signed(2892422, 24), to_signed(2899037, 24), to_signed(2905645, 24), to_signed(2912246, 24), to_signed(2918841, 24), to_signed(2925428, 24), to_signed(2932009, 24), to_signed(2938583, 24), to_signed(2945149, 24), to_signed(2951709, 24), to_signed(2958262, 24), to_signed(2964808, 24), to_signed(2971347, 24), to_signed(2977879, 24), to_signed(2984404, 24), to_signed(2990922, 24), to_signed(2997433, 24), to_signed(3003937, 24), to_signed(3010434, 24), to_signed(3016924, 24), to_signed(3023406, 24), to_signed(3029882, 24), to_signed(3036350, 24), to_signed(3042812, 24), to_signed(3049266, 24), to_signed(3055713, 24), to_signed(3062152, 24), to_signed(3068585, 24), to_signed(3075010, 24), to_signed(3081428, 24), to_signed(3087839, 24), to_signed(3094243, 24), to_signed(3100639, 24), to_signed(3107028, 24), to_signed(3113410, 24), to_signed(3119784, 24), to_signed(3126151, 24), to_signed(3132511, 24), to_signed(3138863, 24), to_signed(3145208, 24), to_signed(3151545, 24), to_signed(3157875, 24), to_signed(3164198, 24), to_signed(3170513, 24), to_signed(3176821, 24), to_signed(3183121, 24), to_signed(3189414, 24), to_signed(3195699, 24), to_signed(3201977, 24), to_signed(3208247, 24), to_signed(3214510, 24), to_signed(3220765, 24), to_signed(3227013, 24), to_signed(3233253, 24), to_signed(3239485, 24), to_signed(3245710, 24), to_signed(3251927, 24), to_signed(3258136, 24), to_signed(3264338, 24), to_signed(3270532, 24), to_signed(3276718, 24), to_signed(3282897, 24), to_signed(3289068, 24), to_signed(3295231, 24), to_signed(3301387, 24), to_signed(3307534, 24), to_signed(3313674, 24), to_signed(3319806, 24), to_signed(3325930, 24), to_signed(3332047, 24), to_signed(3338156, 24), to_signed(3344256, 24), to_signed(3350349, 24), to_signed(3356434, 24), to_signed(3362511, 24), to_signed(3368580, 24), to_signed(3374642, 24), to_signed(3380695, 24), to_signed(3386740, 24), to_signed(3392778, 24), to_signed(3398807, 24), to_signed(3404829, 24), to_signed(3410842, 24), to_signed(3416847, 24), to_signed(3422845, 24), to_signed(3428834, 24), to_signed(3434815, 24), to_signed(3440788, 24), to_signed(3446753, 24), to_signed(3452710, 24), to_signed(3458659, 24), to_signed(3464600, 24), to_signed(3470532, 24), to_signed(3476457, 24), to_signed(3482373, 24), to_signed(3488281, 24), to_signed(3494181, 24), to_signed(3500072, 24), to_signed(3505955, 24), to_signed(3511831, 24), to_signed(3517697, 24), to_signed(3523556, 24), to_signed(3529406, 24), to_signed(3535248, 24), to_signed(3541082, 24), to_signed(3546907, 24), to_signed(3552724, 24), to_signed(3558532, 24), to_signed(3564333, 24), to_signed(3570124, 24), to_signed(3575908, 24), to_signed(3581683, 24), to_signed(3587449, 24), to_signed(3593207, 24), to_signed(3598957, 24), to_signed(3604698, 24), to_signed(3610431, 24), to_signed(3616155, 24), to_signed(3621871, 24), to_signed(3627578, 24), to_signed(3633277, 24), to_signed(3638967, 24), to_signed(3644648, 24), to_signed(3650321, 24), to_signed(3655986, 24), to_signed(3661641, 24), to_signed(3667289, 24), to_signed(3672927, 24), to_signed(3678557, 24), to_signed(3684178, 24), to_signed(3689791, 24), to_signed(3695395, 24), to_signed(3700990, 24), to_signed(3706576, 24), to_signed(3712154, 24), to_signed(3717723, 24), to_signed(3723283, 24), to_signed(3728835, 24), to_signed(3734377, 24), to_signed(3739911, 24), to_signed(3745437, 24), to_signed(3750953, 24), to_signed(3756460, 24), to_signed(3761959, 24), to_signed(3767449, 24), to_signed(3772930, 24), to_signed(3778402, 24), to_signed(3783865, 24), to_signed(3789319, 24), to_signed(3794765, 24), to_signed(3800201, 24), to_signed(3805629, 24), to_signed(3811047, 24), to_signed(3816457, 24), to_signed(3821857, 24), to_signed(3827249, 24), to_signed(3832631, 24), to_signed(3838005, 24), to_signed(3843369, 24), to_signed(3848725, 24), to_signed(3854071, 24), to_signed(3859409, 24), to_signed(3864737, 24), to_signed(3870056, 24), to_signed(3875366, 24), to_signed(3880667, 24), to_signed(3885959, 24), to_signed(3891242, 24), to_signed(3896515, 24), to_signed(3901780, 24), to_signed(3907035, 24), to_signed(3912281, 24), to_signed(3917517, 24), to_signed(3922745, 24), to_signed(3927963, 24), to_signed(3933172, 24), to_signed(3938372, 24), to_signed(3943563, 24), to_signed(3948744, 24), to_signed(3953916, 24), to_signed(3959079, 24), to_signed(3964232, 24), to_signed(3969376, 24), to_signed(3974511, 24), to_signed(3979636, 24), to_signed(3984752, 24), to_signed(3989859, 24), to_signed(3994956, 24), to_signed(4000044, 24), to_signed(4005122, 24), to_signed(4010191, 24), to_signed(4015251, 24), to_signed(4020301, 24), to_signed(4025342, 24), to_signed(4030373, 24), to_signed(4035394, 24), to_signed(4040407, 24), to_signed(4045409, 24), to_signed(4050402, 24), to_signed(4055386, 24), to_signed(4060360, 24), to_signed(4065325, 24), to_signed(4070280, 24), to_signed(4075225, 24), to_signed(4080161, 24), to_signed(4085087, 24), to_signed(4090004, 24), to_signed(4094911, 24), to_signed(4099808, 24), to_signed(4104696, 24), to_signed(4109574, 24), to_signed(4114442, 24), to_signed(4119301, 24), to_signed(4124149, 24), to_signed(4128989, 24), to_signed(4133818, 24), to_signed(4138638, 24), to_signed(4143448, 24), to_signed(4148249, 24), to_signed(4153039, 24), to_signed(4157820, 24), to_signed(4162591, 24), to_signed(4167352, 24), to_signed(4172104, 24), to_signed(4176845, 24), to_signed(4181577, 24), to_signed(4186299, 24), to_signed(4191011, 24), to_signed(4195713, 24), to_signed(4200406, 24), to_signed(4205088, 24), to_signed(4209761, 24), to_signed(4214423, 24), to_signed(4219076, 24), to_signed(4223719, 24), to_signed(4228352, 24), to_signed(4232975, 24), to_signed(4237588, 24), to_signed(4242191, 24), to_signed(4246784, 24), to_signed(4251367, 24), to_signed(4255940, 24), to_signed(4260503, 24), to_signed(4265056, 24), to_signed(4269599, 24), to_signed(4274131, 24), to_signed(4278654, 24), to_signed(4283167, 24), to_signed(4287670, 24), to_signed(4292162, 24), to_signed(4296645, 24), to_signed(4301117, 24), to_signed(4305579, 24), to_signed(4310032, 24), to_signed(4314474, 24), to_signed(4318905, 24), to_signed(4323327, 24), to_signed(4327739, 24), to_signed(4332140, 24), to_signed(4336531, 24), to_signed(4340912, 24), to_signed(4345283, 24), to_signed(4349643, 24), to_signed(4353993, 24), to_signed(4358333, 24), to_signed(4362663, 24), to_signed(4366983, 24), to_signed(4371292, 24), to_signed(4375591, 24), to_signed(4379879, 24), to_signed(4384158, 24), to_signed(4388426, 24), to_signed(4392683, 24), to_signed(4396931, 24), to_signed(4401168, 24), to_signed(4405394, 24), to_signed(4409611, 24), to_signed(4413817, 24), to_signed(4418012, 24), to_signed(4422197, 24), to_signed(4426372, 24), to_signed(4430536, 24), to_signed(4434690, 24), to_signed(4438833, 24), to_signed(4442966, 24), to_signed(4447089, 24), to_signed(4451201, 24), to_signed(4455303, 24), to_signed(4459394, 24), to_signed(4463474, 24), to_signed(4467544, 24), to_signed(4471604, 24), to_signed(4475653, 24), to_signed(4479692, 24), to_signed(4483720, 24), to_signed(4487737, 24), to_signed(4491744, 24), to_signed(4495740, 24), to_signed(4499726, 24), to_signed(4503701, 24), to_signed(4507666, 24), to_signed(4511620, 24), to_signed(4515563, 24), to_signed(4519496, 24), to_signed(4523418, 24), to_signed(4527329, 24), to_signed(4531230, 24), to_signed(4535120, 24), to_signed(4539000, 24), to_signed(4542868, 24), to_signed(4546727, 24), to_signed(4550574, 24), to_signed(4554411, 24), to_signed(4558237, 24), to_signed(4562052, 24), to_signed(4565856, 24), to_signed(4569650, 24), to_signed(4573433, 24), to_signed(4577205, 24), to_signed(4580967, 24), to_signed(4584717, 24), to_signed(4588457, 24), to_signed(4592186, 24), to_signed(4595905, 24), to_signed(4599612, 24), to_signed(4603309, 24), to_signed(4606995, 24), to_signed(4610670, 24), to_signed(4614334, 24), to_signed(4617987, 24), to_signed(4621629, 24), to_signed(4625261, 24), to_signed(4628882, 24), to_signed(4632491, 24), to_signed(4636090, 24), to_signed(4639678, 24), to_signed(4643255, 24), to_signed(4646821, 24), to_signed(4650376, 24), to_signed(4653921, 24), to_signed(4657454, 24), to_signed(4660976, 24), to_signed(4664488, 24), to_signed(4667988, 24), to_signed(4671477, 24), to_signed(4674956, 24), to_signed(4678423, 24), to_signed(4681879, 24), to_signed(4685325, 24), to_signed(4688759, 24), to_signed(4692182, 24), to_signed(4695595, 24), to_signed(4698996, 24), to_signed(4702386, 24), to_signed(4705765, 24), to_signed(4709133, 24), to_signed(4712490, 24), to_signed(4715836, 24), to_signed(4719171, 24), to_signed(4722494, 24), to_signed(4725807, 24), to_signed(4729108, 24), to_signed(4732399, 24), to_signed(4735678, 24), to_signed(4738946, 24), to_signed(4742203, 24), to_signed(4745448, 24), to_signed(4748683, 24), to_signed(4751906, 24), to_signed(4755118, 24), to_signed(4758319, 24), to_signed(4761509, 24), to_signed(4764688, 24), to_signed(4767855, 24), to_signed(4771011, 24), to_signed(4774156, 24), to_signed(4777290, 24), to_signed(4780412, 24), to_signed(4783524, 24), to_signed(4786624, 24), to_signed(4789712, 24), to_signed(4792790, 24), to_signed(4795856, 24), to_signed(4798911, 24), to_signed(4801954, 24), to_signed(4804986, 24), to_signed(4808007, 24), to_signed(4811017, 24), to_signed(4814015, 24), to_signed(4817002, 24), to_signed(4819978, 24), to_signed(4822942, 24), to_signed(4825895, 24), to_signed(4828837, 24), to_signed(4831767, 24), to_signed(4834686, 24), to_signed(4837594, 24), to_signed(4840490, 24), to_signed(4843374, 24), to_signed(4846248, 24), to_signed(4849110, 24), to_signed(4851960, 24), to_signed(4854799, 24), to_signed(4857627, 24), to_signed(4860443, 24), to_signed(4863248, 24), to_signed(4866041, 24), to_signed(4868823, 24), to_signed(4871594, 24), to_signed(4874353, 24), to_signed(4877100, 24), to_signed(4879836, 24), to_signed(4882561, 24), to_signed(4885274, 24), to_signed(4887976, 24), to_signed(4890666, 24), to_signed(4893344, 24), to_signed(4896011, 24), to_signed(4898667, 24), to_signed(4901311, 24), to_signed(4903943, 24), to_signed(4906564, 24), to_signed(4909174, 24), to_signed(4911771, 24), to_signed(4914358, 24), to_signed(4916932, 24), to_signed(4919496, 24), to_signed(4922047, 24), to_signed(4924587, 24), to_signed(4927116, 24), to_signed(4929632, 24), to_signed(4932138, 24), to_signed(4934631, 24), to_signed(4937113, 24), to_signed(4939583, 24), to_signed(4942042, 24), to_signed(4944489, 24), to_signed(4946925, 24), to_signed(4949349, 24), to_signed(4951761, 24), to_signed(4954161, 24), to_signed(4956550, 24), to_signed(4958928, 24), to_signed(4961293, 24), to_signed(4963647, 24), to_signed(4965989, 24), to_signed(4968320, 24), to_signed(4970639, 24), to_signed(4972946, 24), to_signed(4975241, 24), to_signed(4977525, 24), to_signed(4979797, 24), to_signed(4982057, 24), to_signed(4984306, 24), to_signed(4986542, 24), to_signed(4988768, 24), to_signed(4990981, 24), to_signed(4993183, 24), to_signed(4995372, 24), to_signed(4997551, 24), to_signed(4999717, 24), to_signed(5001872, 24), to_signed(5004014, 24), to_signed(5006145, 24), to_signed(5008265, 24), to_signed(5010372, 24), to_signed(5012468, 24), to_signed(5014552, 24), to_signed(5016624, 24), to_signed(5018684, 24), to_signed(5020733, 24), to_signed(5022769, 24), to_signed(5024794, 24), to_signed(5026807, 24), to_signed(5028808, 24), to_signed(5030798, 24), to_signed(5032775, 24), to_signed(5034741, 24), to_signed(5036695, 24), to_signed(5038637, 24), to_signed(5040567, 24), to_signed(5042485, 24), to_signed(5044392, 24), to_signed(5046286, 24), to_signed(5048169, 24), to_signed(5050039, 24), to_signed(5051898, 24), to_signed(5053745, 24), to_signed(5055581, 24), to_signed(5057404, 24), to_signed(5059215, 24), to_signed(5061014, 24), to_signed(5062802, 24), to_signed(5064578, 24), to_signed(5066341, 24), to_signed(5068093, 24), to_signed(5069833, 24), to_signed(5071561, 24), to_signed(5073277, 24), to_signed(5074981, 24), to_signed(5076673, 24), to_signed(5078353, 24), to_signed(5080021, 24), to_signed(5081677, 24), to_signed(5083322, 24), to_signed(5084954, 24), to_signed(5086574, 24), to_signed(5088183, 24), to_signed(5089779, 24), to_signed(5091363, 24), to_signed(5092936, 24), to_signed(5094496, 24), to_signed(5096045, 24), to_signed(5097581, 24), to_signed(5099106, 24), to_signed(5100618, 24), to_signed(5102119, 24), to_signed(5103607, 24), to_signed(5105084, 24), to_signed(5106548, 24), to_signed(5108001, 24), to_signed(5109441, 24), to_signed(5110870, 24), to_signed(5112286, 24), to_signed(5113690, 24), to_signed(5115083, 24), to_signed(5116463, 24), to_signed(5117831, 24), to_signed(5119187, 24), to_signed(5120531, 24), to_signed(5121864, 24), to_signed(5123184, 24), to_signed(5124492, 24), to_signed(5125788, 24), to_signed(5127071, 24), to_signed(5128343, 24), to_signed(5129603, 24), to_signed(5130851, 24), to_signed(5132086, 24), to_signed(5133310, 24), to_signed(5134521, 24), to_signed(5135721, 24), to_signed(5136908, 24), to_signed(5138083, 24), to_signed(5139246, 24), to_signed(5140397, 24), to_signed(5141536, 24), to_signed(5142663, 24), to_signed(5143778, 24), to_signed(5144880, 24), to_signed(5145971, 24), to_signed(5147049, 24), to_signed(5148115, 24), to_signed(5149169, 24), to_signed(5150212, 24), to_signed(5151241, 24), to_signed(5152259, 24), to_signed(5153265, 24), to_signed(5154258, 24), to_signed(5155240, 24), to_signed(5156209, 24), to_signed(5157166, 24), to_signed(5158111, 24), to_signed(5159044, 24), to_signed(5159965, 24), to_signed(5160874, 24), to_signed(5161770, 24), to_signed(5162654, 24), to_signed(5163527, 24), to_signed(5164387, 24), to_signed(5165235, 24), to_signed(5166070, 24), to_signed(5166894, 24), to_signed(5167705, 24), to_signed(5168504, 24), to_signed(5169292, 24), to_signed(5170066, 24), to_signed(5170829, 24), to_signed(5171580, 24), to_signed(5172318, 24), to_signed(5173044, 24), to_signed(5173758, 24), to_signed(5174460, 24), to_signed(5175150, 24), to_signed(5175828, 24), to_signed(5176493, 24), to_signed(5177146, 24), to_signed(5177787, 24), to_signed(5178416, 24), to_signed(5179033, 24), to_signed(5179637, 24), to_signed(5180229, 24), to_signed(5180809, 24), to_signed(5181377, 24), to_signed(5181933, 24), to_signed(5182476, 24), to_signed(5183008, 24), to_signed(5183527, 24), to_signed(5184034, 24), to_signed(5184528, 24), to_signed(5185011, 24), to_signed(5185481, 24), to_signed(5185939, 24), to_signed(5186385, 24), to_signed(5186819, 24), to_signed(5187240, 24), to_signed(5187650, 24), to_signed(5188047, 24), to_signed(5188432, 24), to_signed(5188804, 24), to_signed(5189165, 24), to_signed(5189513, 24), to_signed(5189849, 24), to_signed(5190173, 24), to_signed(5190484, 24), to_signed(5190784, 24), to_signed(5191071, 24), to_signed(5191346, 24), to_signed(5191609, 24), to_signed(5191859, 24), to_signed(5192097, 24), to_signed(5192324, 24), to_signed(5192537, 24), to_signed(5192739, 24), to_signed(5192929, 24), to_signed(5193106, 24), to_signed(5193271, 24), to_signed(5193423, 24), to_signed(5193564, 24), to_signed(5193692, 24), to_signed(5193808, 24), to_signed(5193912, 24), to_signed(5194004, 24), to_signed(5194083, 24), to_signed(5194151, 24), to_signed(5194206, 24), to_signed(5194248, 24), to_signed(5194279, 24), to_signed(5194297, 24), to_signed(5194304, 24), to_signed(5194297, 24), to_signed(5194279, 24), to_signed(5194248, 24), to_signed(5194206, 24), to_signed(5194151, 24), to_signed(5194083, 24), to_signed(5194004, 24), to_signed(5193912, 24), to_signed(5193808, 24), to_signed(5193692, 24), to_signed(5193564, 24), to_signed(5193423, 24), to_signed(5193271, 24), to_signed(5193106, 24), to_signed(5192929, 24), to_signed(5192739, 24), to_signed(5192537, 24), to_signed(5192324, 24), to_signed(5192097, 24), to_signed(5191859, 24), to_signed(5191609, 24), to_signed(5191346, 24), to_signed(5191071, 24), to_signed(5190784, 24), to_signed(5190484, 24), to_signed(5190173, 24), to_signed(5189849, 24), to_signed(5189513, 24), to_signed(5189165, 24), to_signed(5188804, 24), to_signed(5188432, 24), to_signed(5188047, 24), to_signed(5187650, 24), to_signed(5187240, 24), to_signed(5186819, 24), to_signed(5186385, 24), to_signed(5185939, 24), to_signed(5185481, 24), to_signed(5185011, 24), to_signed(5184528, 24), to_signed(5184034, 24), to_signed(5183527, 24), to_signed(5183008, 24), to_signed(5182476, 24), to_signed(5181933, 24), to_signed(5181377, 24), to_signed(5180809, 24), to_signed(5180229, 24), to_signed(5179637, 24), to_signed(5179033, 24), to_signed(5178416, 24), to_signed(5177787, 24), to_signed(5177146, 24), to_signed(5176493, 24), to_signed(5175828, 24), to_signed(5175150, 24), to_signed(5174460, 24), to_signed(5173758, 24), to_signed(5173044, 24), to_signed(5172318, 24), to_signed(5171580, 24), to_signed(5170829, 24), to_signed(5170066, 24), to_signed(5169292, 24), to_signed(5168504, 24), to_signed(5167705, 24), to_signed(5166894, 24), to_signed(5166070, 24), to_signed(5165235, 24), to_signed(5164387, 24), to_signed(5163527, 24), to_signed(5162654, 24), to_signed(5161770, 24), to_signed(5160874, 24), to_signed(5159965, 24), to_signed(5159044, 24), to_signed(5158111, 24), to_signed(5157166, 24), to_signed(5156209, 24), to_signed(5155240, 24), to_signed(5154258, 24), to_signed(5153265, 24), to_signed(5152259, 24), to_signed(5151241, 24), to_signed(5150212, 24), to_signed(5149169, 24), to_signed(5148115, 24), to_signed(5147049, 24), to_signed(5145971, 24), to_signed(5144880, 24), to_signed(5143778, 24), to_signed(5142663, 24), to_signed(5141536, 24), to_signed(5140397, 24), to_signed(5139246, 24), to_signed(5138083, 24), to_signed(5136908, 24), to_signed(5135721, 24), to_signed(5134521, 24), to_signed(5133310, 24), to_signed(5132086, 24), to_signed(5130851, 24), to_signed(5129603, 24), to_signed(5128343, 24), to_signed(5127071, 24), to_signed(5125788, 24), to_signed(5124492, 24), to_signed(5123184, 24), to_signed(5121864, 24), to_signed(5120531, 24), to_signed(5119187, 24), to_signed(5117831, 24), to_signed(5116463, 24), to_signed(5115083, 24), to_signed(5113690, 24), to_signed(5112286, 24), to_signed(5110870, 24), to_signed(5109441, 24), to_signed(5108001, 24), to_signed(5106548, 24), to_signed(5105084, 24), to_signed(5103607, 24), to_signed(5102119, 24), to_signed(5100618, 24), to_signed(5099106, 24), to_signed(5097581, 24), to_signed(5096045, 24), to_signed(5094496, 24), to_signed(5092936, 24), to_signed(5091363, 24), to_signed(5089779, 24), to_signed(5088183, 24), to_signed(5086574, 24), to_signed(5084954, 24), to_signed(5083322, 24), to_signed(5081677, 24), to_signed(5080021, 24), to_signed(5078353, 24), to_signed(5076673, 24), to_signed(5074981, 24), to_signed(5073277, 24), to_signed(5071561, 24), to_signed(5069833, 24), to_signed(5068093, 24), to_signed(5066341, 24), to_signed(5064578, 24), to_signed(5062802, 24), to_signed(5061014, 24), to_signed(5059215, 24), to_signed(5057404, 24), to_signed(5055581, 24), to_signed(5053745, 24), to_signed(5051898, 24), to_signed(5050039, 24), to_signed(5048169, 24), to_signed(5046286, 24), to_signed(5044392, 24), to_signed(5042485, 24), to_signed(5040567, 24), to_signed(5038637, 24), to_signed(5036695, 24), to_signed(5034741, 24), to_signed(5032775, 24), to_signed(5030798, 24), to_signed(5028808, 24), to_signed(5026807, 24), to_signed(5024794, 24), to_signed(5022769, 24), to_signed(5020733, 24), to_signed(5018684, 24), to_signed(5016624, 24), to_signed(5014552, 24), to_signed(5012468, 24), to_signed(5010372, 24), to_signed(5008265, 24), to_signed(5006145, 24), to_signed(5004014, 24), to_signed(5001872, 24), to_signed(4999717, 24), to_signed(4997551, 24), to_signed(4995372, 24), to_signed(4993183, 24), to_signed(4990981, 24), to_signed(4988768, 24), to_signed(4986542, 24), to_signed(4984306, 24), to_signed(4982057, 24), to_signed(4979797, 24), to_signed(4977525, 24), to_signed(4975241, 24), to_signed(4972946, 24), to_signed(4970639, 24), to_signed(4968320, 24), to_signed(4965989, 24), to_signed(4963647, 24), to_signed(4961293, 24), to_signed(4958928, 24), to_signed(4956550, 24), to_signed(4954161, 24), to_signed(4951761, 24), to_signed(4949349, 24), to_signed(4946925, 24), to_signed(4944489, 24), to_signed(4942042, 24), to_signed(4939583, 24), to_signed(4937113, 24), to_signed(4934631, 24), to_signed(4932138, 24), to_signed(4929632, 24), to_signed(4927116, 24), to_signed(4924587, 24), to_signed(4922047, 24), to_signed(4919496, 24), to_signed(4916932, 24), to_signed(4914358, 24), to_signed(4911771, 24), to_signed(4909174, 24), to_signed(4906564, 24), to_signed(4903943, 24), to_signed(4901311, 24), to_signed(4898667, 24), to_signed(4896011, 24), to_signed(4893344, 24), to_signed(4890666, 24), to_signed(4887976, 24), to_signed(4885274, 24), to_signed(4882561, 24), to_signed(4879836, 24), to_signed(4877100, 24), to_signed(4874353, 24), to_signed(4871594, 24), to_signed(4868823, 24), to_signed(4866041, 24), to_signed(4863248, 24), to_signed(4860443, 24), to_signed(4857627, 24), to_signed(4854799, 24), to_signed(4851960, 24), to_signed(4849110, 24), to_signed(4846248, 24), to_signed(4843374, 24), to_signed(4840490, 24), to_signed(4837594, 24), to_signed(4834686, 24), to_signed(4831767, 24), to_signed(4828837, 24), to_signed(4825895, 24), to_signed(4822942, 24), to_signed(4819978, 24), to_signed(4817002, 24), to_signed(4814015, 24), to_signed(4811017, 24), to_signed(4808007, 24), to_signed(4804986, 24), to_signed(4801954, 24), to_signed(4798911, 24), to_signed(4795856, 24), to_signed(4792790, 24), to_signed(4789712, 24), to_signed(4786624, 24), to_signed(4783524, 24), to_signed(4780412, 24), to_signed(4777290, 24), to_signed(4774156, 24), to_signed(4771011, 24), to_signed(4767855, 24), to_signed(4764688, 24), to_signed(4761509, 24), to_signed(4758319, 24), to_signed(4755118, 24), to_signed(4751906, 24), to_signed(4748683, 24), to_signed(4745448, 24), to_signed(4742203, 24), to_signed(4738946, 24), to_signed(4735678, 24), to_signed(4732399, 24), to_signed(4729108, 24), to_signed(4725807, 24), to_signed(4722494, 24), to_signed(4719171, 24), to_signed(4715836, 24), to_signed(4712490, 24), to_signed(4709133, 24), to_signed(4705765, 24), to_signed(4702386, 24), to_signed(4698996, 24), to_signed(4695595, 24), to_signed(4692182, 24), to_signed(4688759, 24), to_signed(4685325, 24), to_signed(4681879, 24), to_signed(4678423, 24), to_signed(4674956, 24), to_signed(4671477, 24), to_signed(4667988, 24), to_signed(4664488, 24), to_signed(4660976, 24), to_signed(4657454, 24), to_signed(4653921, 24), to_signed(4650376, 24), to_signed(4646821, 24), to_signed(4643255, 24), to_signed(4639678, 24), to_signed(4636090, 24), to_signed(4632491, 24), to_signed(4628882, 24), to_signed(4625261, 24), to_signed(4621629, 24), to_signed(4617987, 24), to_signed(4614334, 24), to_signed(4610670, 24), to_signed(4606995, 24), to_signed(4603309, 24), to_signed(4599612, 24), to_signed(4595905, 24), to_signed(4592186, 24), to_signed(4588457, 24), to_signed(4584717, 24), to_signed(4580967, 24), to_signed(4577205, 24), to_signed(4573433, 24), to_signed(4569650, 24), to_signed(4565856, 24), to_signed(4562052, 24), to_signed(4558237, 24), to_signed(4554411, 24), to_signed(4550574, 24), to_signed(4546727, 24), to_signed(4542868, 24), to_signed(4539000, 24), to_signed(4535120, 24), to_signed(4531230, 24), to_signed(4527329, 24), to_signed(4523418, 24), to_signed(4519496, 24), to_signed(4515563, 24), to_signed(4511620, 24), to_signed(4507666, 24), to_signed(4503701, 24), to_signed(4499726, 24), to_signed(4495740, 24), to_signed(4491744, 24), to_signed(4487737, 24), to_signed(4483720, 24), to_signed(4479692, 24), to_signed(4475653, 24), to_signed(4471604, 24), to_signed(4467544, 24), to_signed(4463474, 24), to_signed(4459394, 24), to_signed(4455303, 24), to_signed(4451201, 24), to_signed(4447089, 24), to_signed(4442966, 24), to_signed(4438833, 24), to_signed(4434690, 24), to_signed(4430536, 24), to_signed(4426372, 24), to_signed(4422197, 24), to_signed(4418012, 24), to_signed(4413817, 24), to_signed(4409611, 24), to_signed(4405394, 24), to_signed(4401168, 24), to_signed(4396931, 24), to_signed(4392683, 24), to_signed(4388426, 24), to_signed(4384158, 24), to_signed(4379879, 24), to_signed(4375591, 24), to_signed(4371292, 24), to_signed(4366983, 24), to_signed(4362663, 24), to_signed(4358333, 24), to_signed(4353993, 24), to_signed(4349643, 24), to_signed(4345283, 24), to_signed(4340912, 24), to_signed(4336531, 24), to_signed(4332140, 24), to_signed(4327739, 24), to_signed(4323327, 24), to_signed(4318905, 24), to_signed(4314474, 24), to_signed(4310032, 24), to_signed(4305579, 24), to_signed(4301117, 24), to_signed(4296645, 24), to_signed(4292162, 24), to_signed(4287670, 24), to_signed(4283167, 24), to_signed(4278654, 24), to_signed(4274131, 24), to_signed(4269599, 24), to_signed(4265056, 24), to_signed(4260503, 24), to_signed(4255940, 24), to_signed(4251367, 24), to_signed(4246784, 24), to_signed(4242191, 24), to_signed(4237588, 24), to_signed(4232975, 24), to_signed(4228352, 24), to_signed(4223719, 24), to_signed(4219076, 24), to_signed(4214423, 24), to_signed(4209761, 24), to_signed(4205088, 24), to_signed(4200406, 24), to_signed(4195713, 24), to_signed(4191011, 24), to_signed(4186299, 24), to_signed(4181577, 24), to_signed(4176845, 24), to_signed(4172104, 24), to_signed(4167352, 24), to_signed(4162591, 24), to_signed(4157820, 24), to_signed(4153039, 24), to_signed(4148249, 24), to_signed(4143448, 24), to_signed(4138638, 24), to_signed(4133818, 24), to_signed(4128989, 24), to_signed(4124149, 24), to_signed(4119301, 24), to_signed(4114442, 24), to_signed(4109574, 24), to_signed(4104696, 24), to_signed(4099808, 24), to_signed(4094911, 24), to_signed(4090004, 24), to_signed(4085087, 24), to_signed(4080161, 24), to_signed(4075225, 24), to_signed(4070280, 24), to_signed(4065325, 24), to_signed(4060360, 24), to_signed(4055386, 24), to_signed(4050402, 24), to_signed(4045409, 24), to_signed(4040407, 24), to_signed(4035394, 24), to_signed(4030373, 24), to_signed(4025342, 24), to_signed(4020301, 24), to_signed(4015251, 24), to_signed(4010191, 24), to_signed(4005122, 24), to_signed(4000044, 24), to_signed(3994956, 24), to_signed(3989859, 24), to_signed(3984752, 24), to_signed(3979636, 24), to_signed(3974511, 24), to_signed(3969376, 24), to_signed(3964232, 24), to_signed(3959079, 24), to_signed(3953916, 24), to_signed(3948744, 24), to_signed(3943563, 24), to_signed(3938372, 24), to_signed(3933172, 24), to_signed(3927963, 24), to_signed(3922745, 24), to_signed(3917517, 24), to_signed(3912281, 24), to_signed(3907035, 24), to_signed(3901780, 24), to_signed(3896515, 24), to_signed(3891242, 24), to_signed(3885959, 24), to_signed(3880667, 24), to_signed(3875366, 24), to_signed(3870056, 24), to_signed(3864737, 24), to_signed(3859409, 24), to_signed(3854071, 24), to_signed(3848725, 24), to_signed(3843369, 24), to_signed(3838005, 24), to_signed(3832631, 24), to_signed(3827249, 24), to_signed(3821857, 24), to_signed(3816457, 24), to_signed(3811047, 24), to_signed(3805629, 24), to_signed(3800201, 24), to_signed(3794765, 24), to_signed(3789319, 24), to_signed(3783865, 24), to_signed(3778402, 24), to_signed(3772930, 24), to_signed(3767449, 24), to_signed(3761959, 24), to_signed(3756460, 24), to_signed(3750953, 24), to_signed(3745437, 24), to_signed(3739911, 24), to_signed(3734377, 24), to_signed(3728835, 24), to_signed(3723283, 24), to_signed(3717723, 24), to_signed(3712154, 24), to_signed(3706576, 24), to_signed(3700990, 24), to_signed(3695395, 24), to_signed(3689791, 24), to_signed(3684178, 24), to_signed(3678557, 24), to_signed(3672927, 24), to_signed(3667289, 24), to_signed(3661641, 24), to_signed(3655986, 24), to_signed(3650321, 24), to_signed(3644648, 24), to_signed(3638967, 24), to_signed(3633277, 24), to_signed(3627578, 24), to_signed(3621871, 24), to_signed(3616155, 24), to_signed(3610431, 24), to_signed(3604698, 24), to_signed(3598957, 24), to_signed(3593207, 24), to_signed(3587449, 24), to_signed(3581683, 24), to_signed(3575908, 24), to_signed(3570124, 24), to_signed(3564333, 24), to_signed(3558532, 24), to_signed(3552724, 24), to_signed(3546907, 24), to_signed(3541082, 24), to_signed(3535248, 24), to_signed(3529406, 24), to_signed(3523556, 24), to_signed(3517697, 24), to_signed(3511831, 24), to_signed(3505955, 24), to_signed(3500072, 24), to_signed(3494181, 24), to_signed(3488281, 24), to_signed(3482373, 24), to_signed(3476457, 24), to_signed(3470532, 24), to_signed(3464600, 24), to_signed(3458659, 24), to_signed(3452710, 24), to_signed(3446753, 24), to_signed(3440788, 24), to_signed(3434815, 24), to_signed(3428834, 24), to_signed(3422845, 24), to_signed(3416847, 24), to_signed(3410842, 24), to_signed(3404829, 24), to_signed(3398807, 24), to_signed(3392778, 24), to_signed(3386740, 24), to_signed(3380695, 24), to_signed(3374642, 24), to_signed(3368580, 24), to_signed(3362511, 24), to_signed(3356434, 24), to_signed(3350349, 24), to_signed(3344256, 24), to_signed(3338156, 24), to_signed(3332047, 24), to_signed(3325930, 24), to_signed(3319806, 24), to_signed(3313674, 24), to_signed(3307534, 24), to_signed(3301387, 24), to_signed(3295231, 24), to_signed(3289068, 24), to_signed(3282897, 24), to_signed(3276718, 24), to_signed(3270532, 24), to_signed(3264338, 24), to_signed(3258136, 24), to_signed(3251927, 24), to_signed(3245710, 24), to_signed(3239485, 24), to_signed(3233253, 24), to_signed(3227013, 24), to_signed(3220765, 24), to_signed(3214510, 24), to_signed(3208247, 24), to_signed(3201977, 24), to_signed(3195699, 24), to_signed(3189414, 24), to_signed(3183121, 24), to_signed(3176821, 24), to_signed(3170513, 24), to_signed(3164198, 24), to_signed(3157875, 24), to_signed(3151545, 24), to_signed(3145208, 24), to_signed(3138863, 24), to_signed(3132511, 24), to_signed(3126151, 24), to_signed(3119784, 24), to_signed(3113410, 24), to_signed(3107028, 24), to_signed(3100639, 24), to_signed(3094243, 24), to_signed(3087839, 24), to_signed(3081428, 24), to_signed(3075010, 24), to_signed(3068585, 24), to_signed(3062152, 24), to_signed(3055713, 24), to_signed(3049266, 24), to_signed(3042812, 24), to_signed(3036350, 24), to_signed(3029882, 24), to_signed(3023406, 24), to_signed(3016924, 24), to_signed(3010434, 24), to_signed(3003937, 24), to_signed(2997433, 24), to_signed(2990922, 24), to_signed(2984404, 24), to_signed(2977879, 24), to_signed(2971347, 24), to_signed(2964808, 24), to_signed(2958262, 24), to_signed(2951709, 24), to_signed(2945149, 24), to_signed(2938583, 24), to_signed(2932009, 24), to_signed(2925428, 24), to_signed(2918841, 24), to_signed(2912246, 24), to_signed(2905645, 24), to_signed(2899037, 24), to_signed(2892422, 24), to_signed(2885800, 24), to_signed(2879172, 24), to_signed(2872536, 24), to_signed(2865894, 24), to_signed(2859246, 24), to_signed(2852590, 24), to_signed(2845928, 24), to_signed(2839259, 24), to_signed(2832583, 24), to_signed(2825901, 24), to_signed(2819212, 24), to_signed(2812517, 24), to_signed(2805814, 24), to_signed(2799106, 24), to_signed(2792390, 24), to_signed(2785668, 24), to_signed(2778940, 24), to_signed(2772205, 24), to_signed(2765463, 24), to_signed(2758715, 24), to_signed(2751961, 24), to_signed(2745200, 24), to_signed(2738432, 24), to_signed(2731658, 24), to_signed(2724878, 24), to_signed(2718091, 24), to_signed(2711298, 24), to_signed(2704498, 24), to_signed(2697692, 24), to_signed(2690880, 24), to_signed(2684062, 24), to_signed(2677237, 24), to_signed(2670405, 24), to_signed(2663568, 24), to_signed(2656724, 24), to_signed(2649874, 24), to_signed(2643018, 24), to_signed(2636155, 24), to_signed(2629287, 24), to_signed(2622412, 24), to_signed(2615531, 24), to_signed(2608644, 24), to_signed(2601750, 24), to_signed(2594851, 24), to_signed(2587945, 24), to_signed(2581034, 24), to_signed(2574116, 24), to_signed(2567192, 24), to_signed(2560263, 24), to_signed(2553327, 24), to_signed(2546385, 24), to_signed(2539437, 24), to_signed(2532483, 24), to_signed(2525523, 24), to_signed(2518558, 24), to_signed(2511586, 24), to_signed(2504609, 24), to_signed(2497625, 24), to_signed(2490636, 24), to_signed(2483641, 24), to_signed(2476640, 24), to_signed(2469633, 24), to_signed(2462620, 24), to_signed(2455602, 24), to_signed(2448577, 24), to_signed(2441547, 24), to_signed(2434512, 24), to_signed(2427470, 24), to_signed(2420423, 24), to_signed(2413370, 24), to_signed(2406312, 24), to_signed(2399247, 24), to_signed(2392178, 24), to_signed(2385102, 24), to_signed(2378021, 24), to_signed(2370934, 24), to_signed(2363842, 24), to_signed(2356744, 24), to_signed(2349641, 24), to_signed(2342532, 24), to_signed(2335417, 24), to_signed(2328298, 24), to_signed(2321172, 24), to_signed(2314041, 24), to_signed(2306905, 24), to_signed(2299763, 24), to_signed(2292616, 24), to_signed(2285464, 24), to_signed(2278306, 24), to_signed(2271142, 24), to_signed(2263974, 24), to_signed(2256800, 24), to_signed(2249620, 24), to_signed(2242436, 24), to_signed(2235246, 24), to_signed(2228051, 24), to_signed(2220851, 24), to_signed(2213645, 24), to_signed(2206434, 24), to_signed(2199218, 24), to_signed(2191997, 24), to_signed(2184771, 24), to_signed(2177539, 24), to_signed(2170303, 24), to_signed(2163061, 24), to_signed(2155814, 24), to_signed(2148563, 24), to_signed(2141306, 24), to_signed(2134044, 24), to_signed(2126777, 24), to_signed(2119505, 24), to_signed(2112228, 24), to_signed(2104946, 24), to_signed(2097659, 24), to_signed(2090367, 24), to_signed(2083071, 24), to_signed(2075769, 24), to_signed(2068463, 24), to_signed(2061151, 24), to_signed(2053835, 24), to_signed(2046514, 24), to_signed(2039188, 24), to_signed(2031857, 24), to_signed(2024522, 24), to_signed(2017182, 24), to_signed(2009837, 24), to_signed(2002487, 24), to_signed(1995133, 24), to_signed(1987774, 24), to_signed(1980410, 24), to_signed(1973041, 24), to_signed(1965668, 24), to_signed(1958291, 24), to_signed(1950908, 24), to_signed(1943521, 24), to_signed(1936130, 24), to_signed(1928734, 24), to_signed(1921333, 24), to_signed(1913928, 24), to_signed(1906519, 24), to_signed(1899105, 24), to_signed(1891686, 24), to_signed(1884263, 24), to_signed(1876836, 24), to_signed(1869404, 24), to_signed(1861967, 24), to_signed(1854527, 24), to_signed(1847082, 24), to_signed(1839633, 24), to_signed(1832179, 24), to_signed(1824721, 24), to_signed(1817259, 24), to_signed(1809792, 24), to_signed(1802321, 24), to_signed(1794846, 24), to_signed(1787367, 24), to_signed(1779883, 24), to_signed(1772396, 24), to_signed(1764904, 24), to_signed(1757408, 24), to_signed(1749908, 24), to_signed(1742404, 24), to_signed(1734895, 24), to_signed(1727383, 24), to_signed(1719866, 24), to_signed(1712346, 24), to_signed(1704821, 24), to_signed(1697293, 24), to_signed(1689760, 24), to_signed(1682224, 24), to_signed(1674683, 24), to_signed(1667139, 24), to_signed(1659590, 24), to_signed(1652038, 24), to_signed(1644482, 24), to_signed(1636922, 24), to_signed(1629358, 24), to_signed(1621790, 24), to_signed(1614219, 24), to_signed(1606643, 24), to_signed(1599064, 24), to_signed(1591481, 24), to_signed(1583895, 24), to_signed(1576304, 24), to_signed(1568710, 24), to_signed(1561112, 24), to_signed(1553511, 24), to_signed(1545906, 24), to_signed(1538297, 24), to_signed(1530685, 24), to_signed(1523069, 24), to_signed(1515449, 24), to_signed(1507826, 24), to_signed(1500200, 24), to_signed(1492570, 24), to_signed(1484936, 24), to_signed(1477299, 24), to_signed(1469658, 24), to_signed(1462014, 24), to_signed(1454366, 24), to_signed(1446715, 24), to_signed(1439061, 24), to_signed(1431403, 24), to_signed(1423742, 24), to_signed(1416078, 24), to_signed(1408410, 24), to_signed(1400739, 24), to_signed(1393064, 24), to_signed(1385387, 24), to_signed(1377706, 24), to_signed(1370021, 24), to_signed(1362334, 24), to_signed(1354643, 24), to_signed(1346950, 24), to_signed(1339253, 24), to_signed(1331552, 24), to_signed(1323849, 24), to_signed(1316143, 24), to_signed(1308433, 24), to_signed(1300721, 24), to_signed(1293005, 24), to_signed(1285286, 24), to_signed(1277565, 24), to_signed(1269840, 24), to_signed(1262112, 24), to_signed(1254382, 24), to_signed(1246648, 24), to_signed(1238912, 24), to_signed(1231172, 24), to_signed(1223430, 24), to_signed(1215685, 24), to_signed(1207936, 24), to_signed(1200186, 24), to_signed(1192432, 24), to_signed(1184675, 24), to_signed(1176916, 24), to_signed(1169154, 24), to_signed(1161389, 24), to_signed(1153621, 24), to_signed(1145851, 24), to_signed(1138078, 24), to_signed(1130302, 24), to_signed(1122524, 24), to_signed(1114743, 24), to_signed(1106959, 24), to_signed(1099173, 24), to_signed(1091384, 24), to_signed(1083593, 24), to_signed(1075799, 24), to_signed(1068002, 24), to_signed(1060204, 24), to_signed(1052402, 24), to_signed(1044598, 24), to_signed(1036792, 24), to_signed(1028983, 24), to_signed(1021172, 24), to_signed(1013358, 24), to_signed(1005542, 24), to_signed(997723, 24), to_signed(989903, 24), to_signed(982080, 24), to_signed(974254, 24), to_signed(966427, 24), to_signed(958597, 24), to_signed(950764, 24), to_signed(942930, 24), to_signed(935093, 24), to_signed(927254, 24), to_signed(919413, 24), to_signed(911570, 24), to_signed(903725, 24), to_signed(895877, 24), to_signed(888028, 24), to_signed(880176, 24), to_signed(872322, 24), to_signed(864466, 24), to_signed(856608, 24), to_signed(848749, 24), to_signed(840887, 24), to_signed(833023, 24), to_signed(825157, 24), to_signed(817289, 24), to_signed(809420, 24), to_signed(801548, 24), to_signed(793675, 24), to_signed(785799, 24), to_signed(777922, 24), to_signed(770043, 24), to_signed(762162, 24), to_signed(754280, 24), to_signed(746395, 24), to_signed(738509, 24), to_signed(730621, 24), to_signed(722732, 24), to_signed(714840, 24), to_signed(706947, 24), to_signed(699053, 24), to_signed(691156, 24), to_signed(683258, 24), to_signed(675359, 24), to_signed(667458, 24), to_signed(659555, 24), to_signed(651651, 24), to_signed(643745, 24), to_signed(635838, 24), to_signed(627929, 24), to_signed(620019, 24), to_signed(612107, 24), to_signed(604194, 24), to_signed(596279, 24), to_signed(588363, 24), to_signed(580446, 24), to_signed(572527, 24), to_signed(564607, 24), to_signed(556686, 24), to_signed(548763, 24), to_signed(540839, 24), to_signed(532914, 24), to_signed(524987, 24), to_signed(517059, 24), to_signed(509130, 24), to_signed(501200, 24), to_signed(493269, 24), to_signed(485336, 24), to_signed(477403, 24), to_signed(469468, 24), to_signed(461532, 24), to_signed(453595, 24), to_signed(445657, 24), to_signed(437718, 24), to_signed(429778, 24), to_signed(421836, 24), to_signed(413894, 24), to_signed(405951, 24), to_signed(398007, 24), to_signed(390062, 24), to_signed(382116, 24), to_signed(374169, 24), to_signed(366222, 24), to_signed(358273, 24), to_signed(350324, 24), to_signed(342373, 24), to_signed(334422, 24), to_signed(326471, 24), to_signed(318518, 24), to_signed(310565, 24), to_signed(302611, 24), to_signed(294656, 24), to_signed(286700, 24), to_signed(278744, 24), to_signed(270787, 24), to_signed(262830, 24), to_signed(254872, 24), to_signed(246913, 24), to_signed(238954, 24), to_signed(230994, 24), to_signed(223034, 24), to_signed(215073, 24), to_signed(207112, 24), to_signed(199150, 24), to_signed(191187, 24), to_signed(183225, 24), to_signed(175261, 24), to_signed(167298, 24), to_signed(159334, 24), to_signed(151369, 24), to_signed(143405, 24), to_signed(135440, 24), to_signed(127474, 24), to_signed(119508, 24), to_signed(111542, 24), to_signed(103576, 24), to_signed(95610, 24), to_signed(87643, 24), to_signed(79676, 24), to_signed(71709, 24), to_signed(63742, 24), to_signed(55774, 24), to_signed(47807, 24), to_signed(39839, 24), to_signed(31871, 24), to_signed(23903, 24), to_signed(15935, 24), to_signed(7967, 24), to_signed(0, 24), to_signed(-7967, 24), to_signed(-15935, 24), to_signed(-23903, 24), to_signed(-31871, 24), to_signed(-39839, 24), to_signed(-47807, 24), to_signed(-55774, 24), to_signed(-63742, 24), to_signed(-71709, 24), to_signed(-79676, 24), to_signed(-87643, 24), to_signed(-95610, 24), to_signed(-103576, 24), to_signed(-111542, 24), to_signed(-119508, 24), to_signed(-127474, 24), to_signed(-135440, 24), to_signed(-143405, 24), to_signed(-151369, 24), to_signed(-159334, 24), to_signed(-167298, 24), to_signed(-175261, 24), to_signed(-183225, 24), to_signed(-191187, 24), to_signed(-199150, 24), to_signed(-207112, 24), to_signed(-215073, 24), to_signed(-223034, 24), to_signed(-230994, 24), to_signed(-238954, 24), to_signed(-246913, 24), to_signed(-254872, 24), to_signed(-262830, 24), to_signed(-270787, 24), to_signed(-278744, 24), to_signed(-286700, 24), to_signed(-294656, 24), to_signed(-302611, 24), to_signed(-310565, 24), to_signed(-318518, 24), to_signed(-326471, 24), to_signed(-334422, 24), to_signed(-342373, 24), to_signed(-350324, 24), to_signed(-358273, 24), to_signed(-366222, 24), to_signed(-374169, 24), to_signed(-382116, 24), to_signed(-390062, 24), to_signed(-398007, 24), to_signed(-405951, 24), to_signed(-413894, 24), to_signed(-421836, 24), to_signed(-429778, 24), to_signed(-437718, 24), to_signed(-445657, 24), to_signed(-453595, 24), to_signed(-461532, 24), to_signed(-469468, 24), to_signed(-477403, 24), to_signed(-485336, 24), to_signed(-493269, 24), to_signed(-501200, 24), to_signed(-509130, 24), to_signed(-517059, 24), to_signed(-524987, 24), to_signed(-532914, 24), to_signed(-540839, 24), to_signed(-548763, 24), to_signed(-556686, 24), to_signed(-564607, 24), to_signed(-572527, 24), to_signed(-580446, 24), to_signed(-588363, 24), to_signed(-596279, 24), to_signed(-604194, 24), to_signed(-612107, 24), to_signed(-620019, 24), to_signed(-627929, 24), to_signed(-635838, 24), to_signed(-643745, 24), to_signed(-651651, 24), to_signed(-659555, 24), to_signed(-667458, 24), to_signed(-675359, 24), to_signed(-683258, 24), to_signed(-691156, 24), to_signed(-699053, 24), to_signed(-706947, 24), to_signed(-714840, 24), to_signed(-722732, 24), to_signed(-730621, 24), to_signed(-738509, 24), to_signed(-746395, 24), to_signed(-754280, 24), to_signed(-762162, 24), to_signed(-770043, 24), to_signed(-777922, 24), to_signed(-785799, 24), to_signed(-793675, 24), to_signed(-801548, 24), to_signed(-809420, 24), to_signed(-817289, 24), to_signed(-825157, 24), to_signed(-833023, 24), to_signed(-840887, 24), to_signed(-848749, 24), to_signed(-856608, 24), to_signed(-864466, 24), to_signed(-872322, 24), to_signed(-880176, 24), to_signed(-888028, 24), to_signed(-895877, 24), to_signed(-903725, 24), to_signed(-911570, 24), to_signed(-919413, 24), to_signed(-927254, 24), to_signed(-935093, 24), to_signed(-942930, 24), to_signed(-950764, 24), to_signed(-958597, 24), to_signed(-966427, 24), to_signed(-974254, 24), to_signed(-982080, 24), to_signed(-989903, 24), to_signed(-997723, 24), to_signed(-1005542, 24), to_signed(-1013358, 24), to_signed(-1021172, 24), to_signed(-1028983, 24), to_signed(-1036792, 24), to_signed(-1044598, 24), to_signed(-1052402, 24), to_signed(-1060204, 24), to_signed(-1068002, 24), to_signed(-1075799, 24), to_signed(-1083593, 24), to_signed(-1091384, 24), to_signed(-1099173, 24), to_signed(-1106959, 24), to_signed(-1114743, 24), to_signed(-1122524, 24), to_signed(-1130302, 24), to_signed(-1138078, 24), to_signed(-1145851, 24), to_signed(-1153621, 24), to_signed(-1161389, 24), to_signed(-1169154, 24), to_signed(-1176916, 24), to_signed(-1184675, 24), to_signed(-1192432, 24), to_signed(-1200186, 24), to_signed(-1207936, 24), to_signed(-1215685, 24), to_signed(-1223430, 24), to_signed(-1231172, 24), to_signed(-1238912, 24), to_signed(-1246648, 24), to_signed(-1254382, 24), to_signed(-1262112, 24), to_signed(-1269840, 24), to_signed(-1277565, 24), to_signed(-1285286, 24), to_signed(-1293005, 24), to_signed(-1300721, 24), to_signed(-1308433, 24), to_signed(-1316143, 24), to_signed(-1323849, 24), to_signed(-1331552, 24), to_signed(-1339253, 24), to_signed(-1346950, 24), to_signed(-1354643, 24), to_signed(-1362334, 24), to_signed(-1370021, 24), to_signed(-1377706, 24), to_signed(-1385387, 24), to_signed(-1393064, 24), to_signed(-1400739, 24), to_signed(-1408410, 24), to_signed(-1416078, 24), to_signed(-1423742, 24), to_signed(-1431403, 24), to_signed(-1439061, 24), to_signed(-1446715, 24), to_signed(-1454366, 24), to_signed(-1462014, 24), to_signed(-1469658, 24), to_signed(-1477299, 24), to_signed(-1484936, 24), to_signed(-1492570, 24), to_signed(-1500200, 24), to_signed(-1507826, 24), to_signed(-1515449, 24), to_signed(-1523069, 24), to_signed(-1530685, 24), to_signed(-1538297, 24), to_signed(-1545906, 24), to_signed(-1553511, 24), to_signed(-1561112, 24), to_signed(-1568710, 24), to_signed(-1576304, 24), to_signed(-1583895, 24), to_signed(-1591481, 24), to_signed(-1599064, 24), to_signed(-1606643, 24), to_signed(-1614219, 24), to_signed(-1621790, 24), to_signed(-1629358, 24), to_signed(-1636922, 24), to_signed(-1644482, 24), to_signed(-1652038, 24), to_signed(-1659590, 24), to_signed(-1667139, 24), to_signed(-1674683, 24), to_signed(-1682224, 24), to_signed(-1689760, 24), to_signed(-1697293, 24), to_signed(-1704821, 24), to_signed(-1712346, 24), to_signed(-1719866, 24), to_signed(-1727383, 24), to_signed(-1734895, 24), to_signed(-1742404, 24), to_signed(-1749908, 24), to_signed(-1757408, 24), to_signed(-1764904, 24), to_signed(-1772396, 24), to_signed(-1779883, 24), to_signed(-1787367, 24), to_signed(-1794846, 24), to_signed(-1802321, 24), to_signed(-1809792, 24), to_signed(-1817259, 24), to_signed(-1824721, 24), to_signed(-1832179, 24), to_signed(-1839633, 24), to_signed(-1847082, 24), to_signed(-1854527, 24), to_signed(-1861967, 24), to_signed(-1869404, 24), to_signed(-1876836, 24), to_signed(-1884263, 24), to_signed(-1891686, 24), to_signed(-1899105, 24), to_signed(-1906519, 24), to_signed(-1913928, 24), to_signed(-1921333, 24), to_signed(-1928734, 24), to_signed(-1936130, 24), to_signed(-1943521, 24), to_signed(-1950908, 24), to_signed(-1958291, 24), to_signed(-1965668, 24), to_signed(-1973041, 24), to_signed(-1980410, 24), to_signed(-1987774, 24), to_signed(-1995133, 24), to_signed(-2002487, 24), to_signed(-2009837, 24), to_signed(-2017182, 24), to_signed(-2024522, 24), to_signed(-2031857, 24), to_signed(-2039188, 24), to_signed(-2046514, 24), to_signed(-2053835, 24), to_signed(-2061151, 24), to_signed(-2068463, 24), to_signed(-2075769, 24), to_signed(-2083071, 24), to_signed(-2090367, 24), to_signed(-2097659, 24), to_signed(-2104946, 24), to_signed(-2112228, 24), to_signed(-2119505, 24), to_signed(-2126777, 24), to_signed(-2134044, 24), to_signed(-2141306, 24), to_signed(-2148563, 24), to_signed(-2155814, 24), to_signed(-2163061, 24), to_signed(-2170303, 24), to_signed(-2177539, 24), to_signed(-2184771, 24), to_signed(-2191997, 24), to_signed(-2199218, 24), to_signed(-2206434, 24), to_signed(-2213645, 24), to_signed(-2220851, 24), to_signed(-2228051, 24), to_signed(-2235246, 24), to_signed(-2242436, 24), to_signed(-2249620, 24), to_signed(-2256800, 24), to_signed(-2263974, 24), to_signed(-2271142, 24), to_signed(-2278306, 24), to_signed(-2285464, 24), to_signed(-2292616, 24), to_signed(-2299763, 24), to_signed(-2306905, 24), to_signed(-2314041, 24), to_signed(-2321172, 24), to_signed(-2328298, 24), to_signed(-2335417, 24), to_signed(-2342532, 24), to_signed(-2349641, 24), to_signed(-2356744, 24), to_signed(-2363842, 24), to_signed(-2370934, 24), to_signed(-2378021, 24), to_signed(-2385102, 24), to_signed(-2392178, 24), to_signed(-2399247, 24), to_signed(-2406312, 24), to_signed(-2413370, 24), to_signed(-2420423, 24), to_signed(-2427470, 24), to_signed(-2434512, 24), to_signed(-2441547, 24), to_signed(-2448577, 24), to_signed(-2455602, 24), to_signed(-2462620, 24), to_signed(-2469633, 24), to_signed(-2476640, 24), to_signed(-2483641, 24), to_signed(-2490636, 24), to_signed(-2497625, 24), to_signed(-2504609, 24), to_signed(-2511586, 24), to_signed(-2518558, 24), to_signed(-2525523, 24), to_signed(-2532483, 24), to_signed(-2539437, 24), to_signed(-2546385, 24), to_signed(-2553327, 24), to_signed(-2560263, 24), to_signed(-2567192, 24), to_signed(-2574116, 24), to_signed(-2581034, 24), to_signed(-2587945, 24), to_signed(-2594851, 24), to_signed(-2601750, 24), to_signed(-2608644, 24), to_signed(-2615531, 24), to_signed(-2622412, 24), to_signed(-2629287, 24), to_signed(-2636155, 24), to_signed(-2643018, 24), to_signed(-2649874, 24), to_signed(-2656724, 24), to_signed(-2663568, 24), to_signed(-2670405, 24), to_signed(-2677237, 24), to_signed(-2684062, 24), to_signed(-2690880, 24), to_signed(-2697692, 24), to_signed(-2704498, 24), to_signed(-2711298, 24), to_signed(-2718091, 24), to_signed(-2724878, 24), to_signed(-2731658, 24), to_signed(-2738432, 24), to_signed(-2745200, 24), to_signed(-2751961, 24), to_signed(-2758715, 24), to_signed(-2765463, 24), to_signed(-2772205, 24), to_signed(-2778940, 24), to_signed(-2785668, 24), to_signed(-2792390, 24), to_signed(-2799106, 24), to_signed(-2805814, 24), to_signed(-2812517, 24), to_signed(-2819212, 24), to_signed(-2825901, 24), to_signed(-2832583, 24), to_signed(-2839259, 24), to_signed(-2845928, 24), to_signed(-2852590, 24), to_signed(-2859246, 24), to_signed(-2865894, 24), to_signed(-2872536, 24), to_signed(-2879172, 24), to_signed(-2885800, 24), to_signed(-2892422, 24), to_signed(-2899037, 24), to_signed(-2905645, 24), to_signed(-2912246, 24), to_signed(-2918841, 24), to_signed(-2925428, 24), to_signed(-2932009, 24), to_signed(-2938583, 24), to_signed(-2945149, 24), to_signed(-2951709, 24), to_signed(-2958262, 24), to_signed(-2964808, 24), to_signed(-2971347, 24), to_signed(-2977879, 24), to_signed(-2984404, 24), to_signed(-2990922, 24), to_signed(-2997433, 24), to_signed(-3003937, 24), to_signed(-3010434, 24), to_signed(-3016924, 24), to_signed(-3023406, 24), to_signed(-3029882, 24), to_signed(-3036350, 24), to_signed(-3042812, 24), to_signed(-3049266, 24), to_signed(-3055713, 24), to_signed(-3062152, 24), to_signed(-3068585, 24), to_signed(-3075010, 24), to_signed(-3081428, 24), to_signed(-3087839, 24), to_signed(-3094243, 24), to_signed(-3100639, 24), to_signed(-3107028, 24), to_signed(-3113410, 24), to_signed(-3119784, 24), to_signed(-3126151, 24), to_signed(-3132511, 24), to_signed(-3138863, 24), to_signed(-3145208, 24), to_signed(-3151545, 24), to_signed(-3157875, 24), to_signed(-3164198, 24), to_signed(-3170513, 24), to_signed(-3176821, 24), to_signed(-3183121, 24), to_signed(-3189414, 24), to_signed(-3195699, 24), to_signed(-3201977, 24), to_signed(-3208247, 24), to_signed(-3214510, 24), to_signed(-3220765, 24), to_signed(-3227013, 24), to_signed(-3233253, 24), to_signed(-3239485, 24), to_signed(-3245710, 24), to_signed(-3251927, 24), to_signed(-3258136, 24), to_signed(-3264338, 24), to_signed(-3270532, 24), to_signed(-3276718, 24), to_signed(-3282897, 24), to_signed(-3289068, 24), to_signed(-3295231, 24), to_signed(-3301387, 24), to_signed(-3307534, 24), to_signed(-3313674, 24), to_signed(-3319806, 24), to_signed(-3325930, 24), to_signed(-3332047, 24), to_signed(-3338156, 24), to_signed(-3344256, 24), to_signed(-3350349, 24), to_signed(-3356434, 24), to_signed(-3362511, 24), to_signed(-3368580, 24), to_signed(-3374642, 24), to_signed(-3380695, 24), to_signed(-3386740, 24), to_signed(-3392778, 24), to_signed(-3398807, 24), to_signed(-3404829, 24), to_signed(-3410842, 24), to_signed(-3416847, 24), to_signed(-3422845, 24), to_signed(-3428834, 24), to_signed(-3434815, 24), to_signed(-3440788, 24), to_signed(-3446753, 24), to_signed(-3452710, 24), to_signed(-3458659, 24), to_signed(-3464600, 24), to_signed(-3470532, 24), to_signed(-3476457, 24), to_signed(-3482373, 24), to_signed(-3488281, 24), to_signed(-3494181, 24), to_signed(-3500072, 24), to_signed(-3505955, 24), to_signed(-3511831, 24), to_signed(-3517697, 24), to_signed(-3523556, 24), to_signed(-3529406, 24), to_signed(-3535248, 24), to_signed(-3541082, 24), to_signed(-3546907, 24), to_signed(-3552724, 24), to_signed(-3558532, 24), to_signed(-3564333, 24), to_signed(-3570124, 24), to_signed(-3575908, 24), to_signed(-3581683, 24), to_signed(-3587449, 24), to_signed(-3593207, 24), to_signed(-3598957, 24), to_signed(-3604698, 24), to_signed(-3610431, 24), to_signed(-3616155, 24), to_signed(-3621871, 24), to_signed(-3627578, 24), to_signed(-3633277, 24), to_signed(-3638967, 24), to_signed(-3644648, 24), to_signed(-3650321, 24), to_signed(-3655986, 24), to_signed(-3661641, 24), to_signed(-3667289, 24), to_signed(-3672927, 24), to_signed(-3678557, 24), to_signed(-3684178, 24), to_signed(-3689791, 24), to_signed(-3695395, 24), to_signed(-3700990, 24), to_signed(-3706576, 24), to_signed(-3712154, 24), to_signed(-3717723, 24), to_signed(-3723283, 24), to_signed(-3728835, 24), to_signed(-3734377, 24), to_signed(-3739911, 24), to_signed(-3745437, 24), to_signed(-3750953, 24), to_signed(-3756460, 24), to_signed(-3761959, 24), to_signed(-3767449, 24), to_signed(-3772930, 24), to_signed(-3778402, 24), to_signed(-3783865, 24), to_signed(-3789319, 24), to_signed(-3794765, 24), to_signed(-3800201, 24), to_signed(-3805629, 24), to_signed(-3811047, 24), to_signed(-3816457, 24), to_signed(-3821857, 24), to_signed(-3827249, 24), to_signed(-3832631, 24), to_signed(-3838005, 24), to_signed(-3843369, 24), to_signed(-3848725, 24), to_signed(-3854071, 24), to_signed(-3859409, 24), to_signed(-3864737, 24), to_signed(-3870056, 24), to_signed(-3875366, 24), to_signed(-3880667, 24), to_signed(-3885959, 24), to_signed(-3891242, 24), to_signed(-3896515, 24), to_signed(-3901780, 24), to_signed(-3907035, 24), to_signed(-3912281, 24), to_signed(-3917517, 24), to_signed(-3922745, 24), to_signed(-3927963, 24), to_signed(-3933172, 24), to_signed(-3938372, 24), to_signed(-3943563, 24), to_signed(-3948744, 24), to_signed(-3953916, 24), to_signed(-3959079, 24), to_signed(-3964232, 24), to_signed(-3969376, 24), to_signed(-3974511, 24), to_signed(-3979636, 24), to_signed(-3984752, 24), to_signed(-3989859, 24), to_signed(-3994956, 24), to_signed(-4000044, 24), to_signed(-4005122, 24), to_signed(-4010191, 24), to_signed(-4015251, 24), to_signed(-4020301, 24), to_signed(-4025342, 24), to_signed(-4030373, 24), to_signed(-4035394, 24), to_signed(-4040407, 24), to_signed(-4045409, 24), to_signed(-4050402, 24), to_signed(-4055386, 24), to_signed(-4060360, 24), to_signed(-4065325, 24), to_signed(-4070280, 24), to_signed(-4075225, 24), to_signed(-4080161, 24), to_signed(-4085087, 24), to_signed(-4090004, 24), to_signed(-4094911, 24), to_signed(-4099808, 24), to_signed(-4104696, 24), to_signed(-4109574, 24), to_signed(-4114442, 24), to_signed(-4119301, 24), to_signed(-4124149, 24), to_signed(-4128989, 24), to_signed(-4133818, 24), to_signed(-4138638, 24), to_signed(-4143448, 24), to_signed(-4148249, 24), to_signed(-4153039, 24), to_signed(-4157820, 24), to_signed(-4162591, 24), to_signed(-4167352, 24), to_signed(-4172104, 24), to_signed(-4176845, 24), to_signed(-4181577, 24), to_signed(-4186299, 24), to_signed(-4191011, 24), to_signed(-4195713, 24), to_signed(-4200406, 24), to_signed(-4205088, 24), to_signed(-4209761, 24), to_signed(-4214423, 24), to_signed(-4219076, 24), to_signed(-4223719, 24), to_signed(-4228352, 24), to_signed(-4232975, 24), to_signed(-4237588, 24), to_signed(-4242191, 24), to_signed(-4246784, 24), to_signed(-4251367, 24), to_signed(-4255940, 24), to_signed(-4260503, 24), to_signed(-4265056, 24), to_signed(-4269599, 24), to_signed(-4274131, 24), to_signed(-4278654, 24), to_signed(-4283167, 24), to_signed(-4287670, 24), to_signed(-4292162, 24), to_signed(-4296645, 24), to_signed(-4301117, 24), to_signed(-4305579, 24), to_signed(-4310032, 24), to_signed(-4314474, 24), to_signed(-4318905, 24), to_signed(-4323327, 24), to_signed(-4327739, 24), to_signed(-4332140, 24), to_signed(-4336531, 24), to_signed(-4340912, 24), to_signed(-4345283, 24), to_signed(-4349643, 24), to_signed(-4353993, 24), to_signed(-4358333, 24), to_signed(-4362663, 24), to_signed(-4366983, 24), to_signed(-4371292, 24), to_signed(-4375591, 24), to_signed(-4379879, 24), to_signed(-4384158, 24), to_signed(-4388426, 24), to_signed(-4392683, 24), to_signed(-4396931, 24), to_signed(-4401168, 24), to_signed(-4405394, 24), to_signed(-4409611, 24), to_signed(-4413817, 24), to_signed(-4418012, 24), to_signed(-4422197, 24), to_signed(-4426372, 24), to_signed(-4430536, 24), to_signed(-4434690, 24), to_signed(-4438833, 24), to_signed(-4442966, 24), to_signed(-4447089, 24), to_signed(-4451201, 24), to_signed(-4455303, 24), to_signed(-4459394, 24), to_signed(-4463474, 24), to_signed(-4467544, 24), to_signed(-4471604, 24), to_signed(-4475653, 24), to_signed(-4479692, 24), to_signed(-4483720, 24), to_signed(-4487737, 24), to_signed(-4491744, 24), to_signed(-4495740, 24), to_signed(-4499726, 24), to_signed(-4503701, 24), to_signed(-4507666, 24), to_signed(-4511620, 24), to_signed(-4515563, 24), to_signed(-4519496, 24), to_signed(-4523418, 24), to_signed(-4527329, 24), to_signed(-4531230, 24), to_signed(-4535120, 24), to_signed(-4539000, 24), to_signed(-4542868, 24), to_signed(-4546727, 24), to_signed(-4550574, 24), to_signed(-4554411, 24), to_signed(-4558237, 24), to_signed(-4562052, 24), to_signed(-4565856, 24), to_signed(-4569650, 24), to_signed(-4573433, 24), to_signed(-4577205, 24), to_signed(-4580967, 24), to_signed(-4584717, 24), to_signed(-4588457, 24), to_signed(-4592186, 24), to_signed(-4595905, 24), to_signed(-4599612, 24), to_signed(-4603309, 24), to_signed(-4606995, 24), to_signed(-4610670, 24), to_signed(-4614334, 24), to_signed(-4617987, 24), to_signed(-4621629, 24), to_signed(-4625261, 24), to_signed(-4628882, 24), to_signed(-4632491, 24), to_signed(-4636090, 24), to_signed(-4639678, 24), to_signed(-4643255, 24), to_signed(-4646821, 24), to_signed(-4650376, 24), to_signed(-4653921, 24), to_signed(-4657454, 24), to_signed(-4660976, 24), to_signed(-4664488, 24), to_signed(-4667988, 24), to_signed(-4671477, 24), to_signed(-4674956, 24), to_signed(-4678423, 24), to_signed(-4681879, 24), to_signed(-4685325, 24), to_signed(-4688759, 24), to_signed(-4692182, 24), to_signed(-4695595, 24), to_signed(-4698996, 24), to_signed(-4702386, 24), to_signed(-4705765, 24), to_signed(-4709133, 24), to_signed(-4712490, 24), to_signed(-4715836, 24), to_signed(-4719171, 24), to_signed(-4722494, 24), to_signed(-4725807, 24), to_signed(-4729108, 24), to_signed(-4732399, 24), to_signed(-4735678, 24), to_signed(-4738946, 24), to_signed(-4742203, 24), to_signed(-4745448, 24), to_signed(-4748683, 24), to_signed(-4751906, 24), to_signed(-4755118, 24), to_signed(-4758319, 24), to_signed(-4761509, 24), to_signed(-4764688, 24), to_signed(-4767855, 24), to_signed(-4771011, 24), to_signed(-4774156, 24), to_signed(-4777290, 24), to_signed(-4780412, 24), to_signed(-4783524, 24), to_signed(-4786624, 24), to_signed(-4789712, 24), to_signed(-4792790, 24), to_signed(-4795856, 24), to_signed(-4798911, 24), to_signed(-4801954, 24), to_signed(-4804986, 24), to_signed(-4808007, 24), to_signed(-4811017, 24), to_signed(-4814015, 24), to_signed(-4817002, 24), to_signed(-4819978, 24), to_signed(-4822942, 24), to_signed(-4825895, 24), to_signed(-4828837, 24), to_signed(-4831767, 24), to_signed(-4834686, 24), to_signed(-4837594, 24), to_signed(-4840490, 24), to_signed(-4843374, 24), to_signed(-4846248, 24), to_signed(-4849110, 24), to_signed(-4851960, 24), to_signed(-4854799, 24), to_signed(-4857627, 24), to_signed(-4860443, 24), to_signed(-4863248, 24), to_signed(-4866041, 24), to_signed(-4868823, 24), to_signed(-4871594, 24), to_signed(-4874353, 24), to_signed(-4877100, 24), to_signed(-4879836, 24), to_signed(-4882561, 24), to_signed(-4885274, 24), to_signed(-4887976, 24), to_signed(-4890666, 24), to_signed(-4893344, 24), to_signed(-4896011, 24), to_signed(-4898667, 24), to_signed(-4901311, 24), to_signed(-4903943, 24), to_signed(-4906564, 24), to_signed(-4909174, 24), to_signed(-4911771, 24), to_signed(-4914358, 24), to_signed(-4916932, 24), to_signed(-4919496, 24), to_signed(-4922047, 24), to_signed(-4924587, 24), to_signed(-4927116, 24), to_signed(-4929632, 24), to_signed(-4932138, 24), to_signed(-4934631, 24), to_signed(-4937113, 24), to_signed(-4939583, 24), to_signed(-4942042, 24), to_signed(-4944489, 24), to_signed(-4946925, 24), to_signed(-4949349, 24), to_signed(-4951761, 24), to_signed(-4954161, 24), to_signed(-4956550, 24), to_signed(-4958928, 24), to_signed(-4961293, 24), to_signed(-4963647, 24), to_signed(-4965989, 24), to_signed(-4968320, 24), to_signed(-4970639, 24), to_signed(-4972946, 24), to_signed(-4975241, 24), to_signed(-4977525, 24), to_signed(-4979797, 24), to_signed(-4982057, 24), to_signed(-4984306, 24), to_signed(-4986542, 24), to_signed(-4988768, 24), to_signed(-4990981, 24), to_signed(-4993183, 24), to_signed(-4995372, 24), to_signed(-4997551, 24), to_signed(-4999717, 24), to_signed(-5001872, 24), to_signed(-5004014, 24), to_signed(-5006145, 24), to_signed(-5008265, 24), to_signed(-5010372, 24), to_signed(-5012468, 24), to_signed(-5014552, 24), to_signed(-5016624, 24), to_signed(-5018684, 24), to_signed(-5020733, 24), to_signed(-5022769, 24), to_signed(-5024794, 24), to_signed(-5026807, 24), to_signed(-5028808, 24), to_signed(-5030798, 24), to_signed(-5032775, 24), to_signed(-5034741, 24), to_signed(-5036695, 24), to_signed(-5038637, 24), to_signed(-5040567, 24), to_signed(-5042485, 24), to_signed(-5044392, 24), to_signed(-5046286, 24), to_signed(-5048169, 24), to_signed(-5050039, 24), to_signed(-5051898, 24), to_signed(-5053745, 24), to_signed(-5055581, 24), to_signed(-5057404, 24), to_signed(-5059215, 24), to_signed(-5061014, 24), to_signed(-5062802, 24), to_signed(-5064578, 24), to_signed(-5066341, 24), to_signed(-5068093, 24), to_signed(-5069833, 24), to_signed(-5071561, 24), to_signed(-5073277, 24), to_signed(-5074981, 24), to_signed(-5076673, 24), to_signed(-5078353, 24), to_signed(-5080021, 24), to_signed(-5081677, 24), to_signed(-5083322, 24), to_signed(-5084954, 24), to_signed(-5086574, 24), to_signed(-5088183, 24), to_signed(-5089779, 24), to_signed(-5091363, 24), to_signed(-5092936, 24), to_signed(-5094496, 24), to_signed(-5096045, 24), to_signed(-5097581, 24), to_signed(-5099106, 24), to_signed(-5100618, 24), to_signed(-5102119, 24), to_signed(-5103607, 24), to_signed(-5105084, 24), to_signed(-5106548, 24), to_signed(-5108001, 24), to_signed(-5109441, 24), to_signed(-5110870, 24), to_signed(-5112286, 24), to_signed(-5113690, 24), to_signed(-5115083, 24), to_signed(-5116463, 24), to_signed(-5117831, 24), to_signed(-5119187, 24), to_signed(-5120531, 24), to_signed(-5121864, 24), to_signed(-5123184, 24), to_signed(-5124492, 24), to_signed(-5125788, 24), to_signed(-5127071, 24), to_signed(-5128343, 24), to_signed(-5129603, 24), to_signed(-5130851, 24), to_signed(-5132086, 24), to_signed(-5133310, 24), to_signed(-5134521, 24), to_signed(-5135721, 24), to_signed(-5136908, 24), to_signed(-5138083, 24), to_signed(-5139246, 24), to_signed(-5140397, 24), to_signed(-5141536, 24), to_signed(-5142663, 24), to_signed(-5143778, 24), to_signed(-5144880, 24), to_signed(-5145971, 24), to_signed(-5147049, 24), to_signed(-5148115, 24), to_signed(-5149169, 24), to_signed(-5150212, 24), to_signed(-5151241, 24), to_signed(-5152259, 24), to_signed(-5153265, 24), to_signed(-5154258, 24), to_signed(-5155240, 24), to_signed(-5156209, 24), to_signed(-5157166, 24), to_signed(-5158111, 24), to_signed(-5159044, 24), to_signed(-5159965, 24), to_signed(-5160874, 24), to_signed(-5161770, 24), to_signed(-5162654, 24), to_signed(-5163527, 24), to_signed(-5164387, 24), to_signed(-5165235, 24), to_signed(-5166070, 24), to_signed(-5166894, 24), to_signed(-5167705, 24), to_signed(-5168504, 24), to_signed(-5169292, 24), to_signed(-5170066, 24), to_signed(-5170829, 24), to_signed(-5171580, 24), to_signed(-5172318, 24), to_signed(-5173044, 24), to_signed(-5173758, 24), to_signed(-5174460, 24), to_signed(-5175150, 24), to_signed(-5175828, 24), to_signed(-5176493, 24), to_signed(-5177146, 24), to_signed(-5177787, 24), to_signed(-5178416, 24), to_signed(-5179033, 24), to_signed(-5179637, 24), to_signed(-5180229, 24), to_signed(-5180809, 24), to_signed(-5181377, 24), to_signed(-5181933, 24), to_signed(-5182476, 24), to_signed(-5183008, 24), to_signed(-5183527, 24), to_signed(-5184034, 24), to_signed(-5184528, 24), to_signed(-5185011, 24), to_signed(-5185481, 24), to_signed(-5185939, 24), to_signed(-5186385, 24), to_signed(-5186819, 24), to_signed(-5187240, 24), to_signed(-5187650, 24), to_signed(-5188047, 24), to_signed(-5188432, 24), to_signed(-5188804, 24), to_signed(-5189165, 24), to_signed(-5189513, 24), to_signed(-5189849, 24), to_signed(-5190173, 24), to_signed(-5190484, 24), to_signed(-5190784, 24), to_signed(-5191071, 24), to_signed(-5191346, 24), to_signed(-5191609, 24), to_signed(-5191859, 24), to_signed(-5192097, 24), to_signed(-5192324, 24), to_signed(-5192537, 24), to_signed(-5192739, 24), to_signed(-5192929, 24), to_signed(-5193106, 24), to_signed(-5193271, 24), to_signed(-5193423, 24), to_signed(-5193564, 24), to_signed(-5193692, 24), to_signed(-5193808, 24), to_signed(-5193912, 24), to_signed(-5194004, 24), to_signed(-5194083, 24), to_signed(-5194151, 24), to_signed(-5194206, 24), to_signed(-5194248, 24), to_signed(-5194279, 24), to_signed(-5194297, 24), to_signed(-5194304, 24), to_signed(-5194297, 24), to_signed(-5194279, 24), to_signed(-5194248, 24), to_signed(-5194206, 24), to_signed(-5194151, 24), to_signed(-5194083, 24), to_signed(-5194004, 24), to_signed(-5193912, 24), to_signed(-5193808, 24), to_signed(-5193692, 24), to_signed(-5193564, 24), to_signed(-5193423, 24), to_signed(-5193271, 24), to_signed(-5193106, 24), to_signed(-5192929, 24), to_signed(-5192739, 24), to_signed(-5192537, 24), to_signed(-5192324, 24), to_signed(-5192097, 24), to_signed(-5191859, 24), to_signed(-5191609, 24), to_signed(-5191346, 24), to_signed(-5191071, 24), to_signed(-5190784, 24), to_signed(-5190484, 24), to_signed(-5190173, 24), to_signed(-5189849, 24), to_signed(-5189513, 24), to_signed(-5189165, 24), to_signed(-5188804, 24), to_signed(-5188432, 24), to_signed(-5188047, 24), to_signed(-5187650, 24), to_signed(-5187240, 24), to_signed(-5186819, 24), to_signed(-5186385, 24), to_signed(-5185939, 24), to_signed(-5185481, 24), to_signed(-5185011, 24), to_signed(-5184528, 24), to_signed(-5184034, 24), to_signed(-5183527, 24), to_signed(-5183008, 24), to_signed(-5182476, 24), to_signed(-5181933, 24), to_signed(-5181377, 24), to_signed(-5180809, 24), to_signed(-5180229, 24), to_signed(-5179637, 24), to_signed(-5179033, 24), to_signed(-5178416, 24), to_signed(-5177787, 24), to_signed(-5177146, 24), to_signed(-5176493, 24), to_signed(-5175828, 24), to_signed(-5175150, 24), to_signed(-5174460, 24), to_signed(-5173758, 24), to_signed(-5173044, 24), to_signed(-5172318, 24), to_signed(-5171580, 24), to_signed(-5170829, 24), to_signed(-5170066, 24), to_signed(-5169292, 24), to_signed(-5168504, 24), to_signed(-5167705, 24), to_signed(-5166894, 24), to_signed(-5166070, 24), to_signed(-5165235, 24), to_signed(-5164387, 24), to_signed(-5163527, 24), to_signed(-5162654, 24), to_signed(-5161770, 24), to_signed(-5160874, 24), to_signed(-5159965, 24), to_signed(-5159044, 24), to_signed(-5158111, 24), to_signed(-5157166, 24), to_signed(-5156209, 24), to_signed(-5155240, 24), to_signed(-5154258, 24), to_signed(-5153265, 24), to_signed(-5152259, 24), to_signed(-5151241, 24), to_signed(-5150212, 24), to_signed(-5149169, 24), to_signed(-5148115, 24), to_signed(-5147049, 24), to_signed(-5145971, 24), to_signed(-5144880, 24), to_signed(-5143778, 24), to_signed(-5142663, 24), to_signed(-5141536, 24), to_signed(-5140397, 24), to_signed(-5139246, 24), to_signed(-5138083, 24), to_signed(-5136908, 24), to_signed(-5135721, 24), to_signed(-5134521, 24), to_signed(-5133310, 24), to_signed(-5132086, 24), to_signed(-5130851, 24), to_signed(-5129603, 24), to_signed(-5128343, 24), to_signed(-5127071, 24), to_signed(-5125788, 24), to_signed(-5124492, 24), to_signed(-5123184, 24), to_signed(-5121864, 24), to_signed(-5120531, 24), to_signed(-5119187, 24), to_signed(-5117831, 24), to_signed(-5116463, 24), to_signed(-5115083, 24), to_signed(-5113690, 24), to_signed(-5112286, 24), to_signed(-5110870, 24), to_signed(-5109441, 24), to_signed(-5108001, 24), to_signed(-5106548, 24), to_signed(-5105084, 24), to_signed(-5103607, 24), to_signed(-5102119, 24), to_signed(-5100618, 24), to_signed(-5099106, 24), to_signed(-5097581, 24), to_signed(-5096045, 24), to_signed(-5094496, 24), to_signed(-5092936, 24), to_signed(-5091363, 24), to_signed(-5089779, 24), to_signed(-5088183, 24), to_signed(-5086574, 24), to_signed(-5084954, 24), to_signed(-5083322, 24), to_signed(-5081677, 24), to_signed(-5080021, 24), to_signed(-5078353, 24), to_signed(-5076673, 24), to_signed(-5074981, 24), to_signed(-5073277, 24), to_signed(-5071561, 24), to_signed(-5069833, 24), to_signed(-5068093, 24), to_signed(-5066341, 24), to_signed(-5064578, 24), to_signed(-5062802, 24), to_signed(-5061014, 24), to_signed(-5059215, 24), to_signed(-5057404, 24), to_signed(-5055581, 24), to_signed(-5053745, 24), to_signed(-5051898, 24), to_signed(-5050039, 24), to_signed(-5048169, 24), to_signed(-5046286, 24), to_signed(-5044392, 24), to_signed(-5042485, 24), to_signed(-5040567, 24), to_signed(-5038637, 24), to_signed(-5036695, 24), to_signed(-5034741, 24), to_signed(-5032775, 24), to_signed(-5030798, 24), to_signed(-5028808, 24), to_signed(-5026807, 24), to_signed(-5024794, 24), to_signed(-5022769, 24), to_signed(-5020733, 24), to_signed(-5018684, 24), to_signed(-5016624, 24), to_signed(-5014552, 24), to_signed(-5012468, 24), to_signed(-5010372, 24), to_signed(-5008265, 24), to_signed(-5006145, 24), to_signed(-5004014, 24), to_signed(-5001872, 24), to_signed(-4999717, 24), to_signed(-4997551, 24), to_signed(-4995372, 24), to_signed(-4993183, 24), to_signed(-4990981, 24), to_signed(-4988768, 24), to_signed(-4986542, 24), to_signed(-4984306, 24), to_signed(-4982057, 24), to_signed(-4979797, 24), to_signed(-4977525, 24), to_signed(-4975241, 24), to_signed(-4972946, 24), to_signed(-4970639, 24), to_signed(-4968320, 24), to_signed(-4965989, 24), to_signed(-4963647, 24), to_signed(-4961293, 24), to_signed(-4958928, 24), to_signed(-4956550, 24), to_signed(-4954161, 24), to_signed(-4951761, 24), to_signed(-4949349, 24), to_signed(-4946925, 24), to_signed(-4944489, 24), to_signed(-4942042, 24), to_signed(-4939583, 24), to_signed(-4937113, 24), to_signed(-4934631, 24), to_signed(-4932138, 24), to_signed(-4929632, 24), to_signed(-4927116, 24), to_signed(-4924587, 24), to_signed(-4922047, 24), to_signed(-4919496, 24), to_signed(-4916932, 24), to_signed(-4914358, 24), to_signed(-4911771, 24), to_signed(-4909174, 24), to_signed(-4906564, 24), to_signed(-4903943, 24), to_signed(-4901311, 24), to_signed(-4898667, 24), to_signed(-4896011, 24), to_signed(-4893344, 24), to_signed(-4890666, 24), to_signed(-4887976, 24), to_signed(-4885274, 24), to_signed(-4882561, 24), to_signed(-4879836, 24), to_signed(-4877100, 24), to_signed(-4874353, 24), to_signed(-4871594, 24), to_signed(-4868823, 24), to_signed(-4866041, 24), to_signed(-4863248, 24), to_signed(-4860443, 24), to_signed(-4857627, 24), to_signed(-4854799, 24), to_signed(-4851960, 24), to_signed(-4849110, 24), to_signed(-4846248, 24), to_signed(-4843374, 24), to_signed(-4840490, 24), to_signed(-4837594, 24), to_signed(-4834686, 24), to_signed(-4831767, 24), to_signed(-4828837, 24), to_signed(-4825895, 24), to_signed(-4822942, 24), to_signed(-4819978, 24), to_signed(-4817002, 24), to_signed(-4814015, 24), to_signed(-4811017, 24), to_signed(-4808007, 24), to_signed(-4804986, 24), to_signed(-4801954, 24), to_signed(-4798911, 24), to_signed(-4795856, 24), to_signed(-4792790, 24), to_signed(-4789712, 24), to_signed(-4786624, 24), to_signed(-4783524, 24), to_signed(-4780412, 24), to_signed(-4777290, 24), to_signed(-4774156, 24), to_signed(-4771011, 24), to_signed(-4767855, 24), to_signed(-4764688, 24), to_signed(-4761509, 24), to_signed(-4758319, 24), to_signed(-4755118, 24), to_signed(-4751906, 24), to_signed(-4748683, 24), to_signed(-4745448, 24), to_signed(-4742203, 24), to_signed(-4738946, 24), to_signed(-4735678, 24), to_signed(-4732399, 24), to_signed(-4729108, 24), to_signed(-4725807, 24), to_signed(-4722494, 24), to_signed(-4719171, 24), to_signed(-4715836, 24), to_signed(-4712490, 24), to_signed(-4709133, 24), to_signed(-4705765, 24), to_signed(-4702386, 24), to_signed(-4698996, 24), to_signed(-4695595, 24), to_signed(-4692182, 24), to_signed(-4688759, 24), to_signed(-4685325, 24), to_signed(-4681879, 24), to_signed(-4678423, 24), to_signed(-4674956, 24), to_signed(-4671477, 24), to_signed(-4667988, 24), to_signed(-4664488, 24), to_signed(-4660976, 24), to_signed(-4657454, 24), to_signed(-4653921, 24), to_signed(-4650376, 24), to_signed(-4646821, 24), to_signed(-4643255, 24), to_signed(-4639678, 24), to_signed(-4636090, 24), to_signed(-4632491, 24), to_signed(-4628882, 24), to_signed(-4625261, 24), to_signed(-4621629, 24), to_signed(-4617987, 24), to_signed(-4614334, 24), to_signed(-4610670, 24), to_signed(-4606995, 24), to_signed(-4603309, 24), to_signed(-4599612, 24), to_signed(-4595905, 24), to_signed(-4592186, 24), to_signed(-4588457, 24), to_signed(-4584717, 24), to_signed(-4580967, 24), to_signed(-4577205, 24), to_signed(-4573433, 24), to_signed(-4569650, 24), to_signed(-4565856, 24), to_signed(-4562052, 24), to_signed(-4558237, 24), to_signed(-4554411, 24), to_signed(-4550574, 24), to_signed(-4546727, 24), to_signed(-4542868, 24), to_signed(-4539000, 24), to_signed(-4535120, 24), to_signed(-4531230, 24), to_signed(-4527329, 24), to_signed(-4523418, 24), to_signed(-4519496, 24), to_signed(-4515563, 24), to_signed(-4511620, 24), to_signed(-4507666, 24), to_signed(-4503701, 24), to_signed(-4499726, 24), to_signed(-4495740, 24), to_signed(-4491744, 24), to_signed(-4487737, 24), to_signed(-4483720, 24), to_signed(-4479692, 24), to_signed(-4475653, 24), to_signed(-4471604, 24), to_signed(-4467544, 24), to_signed(-4463474, 24), to_signed(-4459394, 24), to_signed(-4455303, 24), to_signed(-4451201, 24), to_signed(-4447089, 24), to_signed(-4442966, 24), to_signed(-4438833, 24), to_signed(-4434690, 24), to_signed(-4430536, 24), to_signed(-4426372, 24), to_signed(-4422197, 24), to_signed(-4418012, 24), to_signed(-4413817, 24), to_signed(-4409611, 24), to_signed(-4405394, 24), to_signed(-4401168, 24), to_signed(-4396931, 24), to_signed(-4392683, 24), to_signed(-4388426, 24), to_signed(-4384158, 24), to_signed(-4379879, 24), to_signed(-4375591, 24), to_signed(-4371292, 24), to_signed(-4366983, 24), to_signed(-4362663, 24), to_signed(-4358333, 24), to_signed(-4353993, 24), to_signed(-4349643, 24), to_signed(-4345283, 24), to_signed(-4340912, 24), to_signed(-4336531, 24), to_signed(-4332140, 24), to_signed(-4327739, 24), to_signed(-4323327, 24), to_signed(-4318905, 24), to_signed(-4314474, 24), to_signed(-4310032, 24), to_signed(-4305579, 24), to_signed(-4301117, 24), to_signed(-4296645, 24), to_signed(-4292162, 24), to_signed(-4287670, 24), to_signed(-4283167, 24), to_signed(-4278654, 24), to_signed(-4274131, 24), to_signed(-4269599, 24), to_signed(-4265056, 24), to_signed(-4260503, 24), to_signed(-4255940, 24), to_signed(-4251367, 24), to_signed(-4246784, 24), to_signed(-4242191, 24), to_signed(-4237588, 24), to_signed(-4232975, 24), to_signed(-4228352, 24), to_signed(-4223719, 24), to_signed(-4219076, 24), to_signed(-4214423, 24), to_signed(-4209761, 24), to_signed(-4205088, 24), to_signed(-4200406, 24), to_signed(-4195713, 24), to_signed(-4191011, 24), to_signed(-4186299, 24), to_signed(-4181577, 24), to_signed(-4176845, 24), to_signed(-4172104, 24), to_signed(-4167352, 24), to_signed(-4162591, 24), to_signed(-4157820, 24), to_signed(-4153039, 24), to_signed(-4148249, 24), to_signed(-4143448, 24), to_signed(-4138638, 24), to_signed(-4133818, 24), to_signed(-4128989, 24), to_signed(-4124149, 24), to_signed(-4119301, 24), to_signed(-4114442, 24), to_signed(-4109574, 24), to_signed(-4104696, 24), to_signed(-4099808, 24), to_signed(-4094911, 24), to_signed(-4090004, 24), to_signed(-4085087, 24), to_signed(-4080161, 24), to_signed(-4075225, 24), to_signed(-4070280, 24), to_signed(-4065325, 24), to_signed(-4060360, 24), to_signed(-4055386, 24), to_signed(-4050402, 24), to_signed(-4045409, 24), to_signed(-4040407, 24), to_signed(-4035394, 24), to_signed(-4030373, 24), to_signed(-4025342, 24), to_signed(-4020301, 24), to_signed(-4015251, 24), to_signed(-4010191, 24), to_signed(-4005122, 24), to_signed(-4000044, 24), to_signed(-3994956, 24), to_signed(-3989859, 24), to_signed(-3984752, 24), to_signed(-3979636, 24), to_signed(-3974511, 24), to_signed(-3969376, 24), to_signed(-3964232, 24), to_signed(-3959079, 24), to_signed(-3953916, 24), to_signed(-3948744, 24), to_signed(-3943563, 24), to_signed(-3938372, 24), to_signed(-3933172, 24), to_signed(-3927963, 24), to_signed(-3922745, 24), to_signed(-3917517, 24), to_signed(-3912281, 24), to_signed(-3907035, 24), to_signed(-3901780, 24), to_signed(-3896515, 24), to_signed(-3891242, 24), to_signed(-3885959, 24), to_signed(-3880667, 24), to_signed(-3875366, 24), to_signed(-3870056, 24), to_signed(-3864737, 24), to_signed(-3859409, 24), to_signed(-3854071, 24), to_signed(-3848725, 24), to_signed(-3843369, 24), to_signed(-3838005, 24), to_signed(-3832631, 24), to_signed(-3827249, 24), to_signed(-3821857, 24), to_signed(-3816457, 24), to_signed(-3811047, 24), to_signed(-3805629, 24), to_signed(-3800201, 24), to_signed(-3794765, 24), to_signed(-3789319, 24), to_signed(-3783865, 24), to_signed(-3778402, 24), to_signed(-3772930, 24), to_signed(-3767449, 24), to_signed(-3761959, 24), to_signed(-3756460, 24), to_signed(-3750953, 24), to_signed(-3745437, 24), to_signed(-3739911, 24), to_signed(-3734377, 24), to_signed(-3728835, 24), to_signed(-3723283, 24), to_signed(-3717723, 24), to_signed(-3712154, 24), to_signed(-3706576, 24), to_signed(-3700990, 24), to_signed(-3695395, 24), to_signed(-3689791, 24), to_signed(-3684178, 24), to_signed(-3678557, 24), to_signed(-3672927, 24), to_signed(-3667289, 24), to_signed(-3661641, 24), to_signed(-3655986, 24), to_signed(-3650321, 24), to_signed(-3644648, 24), to_signed(-3638967, 24), to_signed(-3633277, 24), to_signed(-3627578, 24), to_signed(-3621871, 24), to_signed(-3616155, 24), to_signed(-3610431, 24), to_signed(-3604698, 24), to_signed(-3598957, 24), to_signed(-3593207, 24), to_signed(-3587449, 24), to_signed(-3581683, 24), to_signed(-3575908, 24), to_signed(-3570124, 24), to_signed(-3564333, 24), to_signed(-3558532, 24), to_signed(-3552724, 24), to_signed(-3546907, 24), to_signed(-3541082, 24), to_signed(-3535248, 24), to_signed(-3529406, 24), to_signed(-3523556, 24), to_signed(-3517697, 24), to_signed(-3511831, 24), to_signed(-3505955, 24), to_signed(-3500072, 24), to_signed(-3494181, 24), to_signed(-3488281, 24), to_signed(-3482373, 24), to_signed(-3476457, 24), to_signed(-3470532, 24), to_signed(-3464600, 24), to_signed(-3458659, 24), to_signed(-3452710, 24), to_signed(-3446753, 24), to_signed(-3440788, 24), to_signed(-3434815, 24), to_signed(-3428834, 24), to_signed(-3422845, 24), to_signed(-3416847, 24), to_signed(-3410842, 24), to_signed(-3404829, 24), to_signed(-3398807, 24), to_signed(-3392778, 24), to_signed(-3386740, 24), to_signed(-3380695, 24), to_signed(-3374642, 24), to_signed(-3368580, 24), to_signed(-3362511, 24), to_signed(-3356434, 24), to_signed(-3350349, 24), to_signed(-3344256, 24), to_signed(-3338156, 24), to_signed(-3332047, 24), to_signed(-3325930, 24), to_signed(-3319806, 24), to_signed(-3313674, 24), to_signed(-3307534, 24), to_signed(-3301387, 24), to_signed(-3295231, 24), to_signed(-3289068, 24), to_signed(-3282897, 24), to_signed(-3276718, 24), to_signed(-3270532, 24), to_signed(-3264338, 24), to_signed(-3258136, 24), to_signed(-3251927, 24), to_signed(-3245710, 24), to_signed(-3239485, 24), to_signed(-3233253, 24), to_signed(-3227013, 24), to_signed(-3220765, 24), to_signed(-3214510, 24), to_signed(-3208247, 24), to_signed(-3201977, 24), to_signed(-3195699, 24), to_signed(-3189414, 24), to_signed(-3183121, 24), to_signed(-3176821, 24), to_signed(-3170513, 24), to_signed(-3164198, 24), to_signed(-3157875, 24), to_signed(-3151545, 24), to_signed(-3145208, 24), to_signed(-3138863, 24), to_signed(-3132511, 24), to_signed(-3126151, 24), to_signed(-3119784, 24), to_signed(-3113410, 24), to_signed(-3107028, 24), to_signed(-3100639, 24), to_signed(-3094243, 24), to_signed(-3087839, 24), to_signed(-3081428, 24), to_signed(-3075010, 24), to_signed(-3068585, 24), to_signed(-3062152, 24), to_signed(-3055713, 24), to_signed(-3049266, 24), to_signed(-3042812, 24), to_signed(-3036350, 24), to_signed(-3029882, 24), to_signed(-3023406, 24), to_signed(-3016924, 24), to_signed(-3010434, 24), to_signed(-3003937, 24), to_signed(-2997433, 24), to_signed(-2990922, 24), to_signed(-2984404, 24), to_signed(-2977879, 24), to_signed(-2971347, 24), to_signed(-2964808, 24), to_signed(-2958262, 24), to_signed(-2951709, 24), to_signed(-2945149, 24), to_signed(-2938583, 24), to_signed(-2932009, 24), to_signed(-2925428, 24), to_signed(-2918841, 24), to_signed(-2912246, 24), to_signed(-2905645, 24), to_signed(-2899037, 24), to_signed(-2892422, 24), to_signed(-2885800, 24), to_signed(-2879172, 24), to_signed(-2872536, 24), to_signed(-2865894, 24), to_signed(-2859246, 24), to_signed(-2852590, 24), to_signed(-2845928, 24), to_signed(-2839259, 24), to_signed(-2832583, 24), to_signed(-2825901, 24), to_signed(-2819212, 24), to_signed(-2812517, 24), to_signed(-2805814, 24), to_signed(-2799106, 24), to_signed(-2792390, 24), to_signed(-2785668, 24), to_signed(-2778940, 24), to_signed(-2772205, 24), to_signed(-2765463, 24), to_signed(-2758715, 24), to_signed(-2751961, 24), to_signed(-2745200, 24), to_signed(-2738432, 24), to_signed(-2731658, 24), to_signed(-2724878, 24), to_signed(-2718091, 24), to_signed(-2711298, 24), to_signed(-2704498, 24), to_signed(-2697692, 24), to_signed(-2690880, 24), to_signed(-2684062, 24), to_signed(-2677237, 24), to_signed(-2670405, 24), to_signed(-2663568, 24), to_signed(-2656724, 24), to_signed(-2649874, 24), to_signed(-2643018, 24), to_signed(-2636155, 24), to_signed(-2629287, 24), to_signed(-2622412, 24), to_signed(-2615531, 24), to_signed(-2608644, 24), to_signed(-2601750, 24), to_signed(-2594851, 24), to_signed(-2587945, 24), to_signed(-2581034, 24), to_signed(-2574116, 24), to_signed(-2567192, 24), to_signed(-2560263, 24), to_signed(-2553327, 24), to_signed(-2546385, 24), to_signed(-2539437, 24), to_signed(-2532483, 24), to_signed(-2525523, 24), to_signed(-2518558, 24), to_signed(-2511586, 24), to_signed(-2504609, 24), to_signed(-2497625, 24), to_signed(-2490636, 24), to_signed(-2483641, 24), to_signed(-2476640, 24), to_signed(-2469633, 24), to_signed(-2462620, 24), to_signed(-2455602, 24), to_signed(-2448577, 24), to_signed(-2441547, 24), to_signed(-2434512, 24), to_signed(-2427470, 24), to_signed(-2420423, 24), to_signed(-2413370, 24), to_signed(-2406312, 24), to_signed(-2399247, 24), to_signed(-2392178, 24), to_signed(-2385102, 24), to_signed(-2378021, 24), to_signed(-2370934, 24), to_signed(-2363842, 24), to_signed(-2356744, 24), to_signed(-2349641, 24), to_signed(-2342532, 24), to_signed(-2335417, 24), to_signed(-2328298, 24), to_signed(-2321172, 24), to_signed(-2314041, 24), to_signed(-2306905, 24), to_signed(-2299763, 24), to_signed(-2292616, 24), to_signed(-2285464, 24), to_signed(-2278306, 24), to_signed(-2271142, 24), to_signed(-2263974, 24), to_signed(-2256800, 24), to_signed(-2249620, 24), to_signed(-2242436, 24), to_signed(-2235246, 24), to_signed(-2228051, 24), to_signed(-2220851, 24), to_signed(-2213645, 24), to_signed(-2206434, 24), to_signed(-2199218, 24), to_signed(-2191997, 24), to_signed(-2184771, 24), to_signed(-2177539, 24), to_signed(-2170303, 24), to_signed(-2163061, 24), to_signed(-2155814, 24), to_signed(-2148563, 24), to_signed(-2141306, 24), to_signed(-2134044, 24), to_signed(-2126777, 24), to_signed(-2119505, 24), to_signed(-2112228, 24), to_signed(-2104946, 24), to_signed(-2097659, 24), to_signed(-2090367, 24), to_signed(-2083071, 24), to_signed(-2075769, 24), to_signed(-2068463, 24), to_signed(-2061151, 24), to_signed(-2053835, 24), to_signed(-2046514, 24), to_signed(-2039188, 24), to_signed(-2031857, 24), to_signed(-2024522, 24), to_signed(-2017182, 24), to_signed(-2009837, 24), to_signed(-2002487, 24), to_signed(-1995133, 24), to_signed(-1987774, 24), to_signed(-1980410, 24), to_signed(-1973041, 24), to_signed(-1965668, 24), to_signed(-1958291, 24), to_signed(-1950908, 24), to_signed(-1943521, 24), to_signed(-1936130, 24), to_signed(-1928734, 24), to_signed(-1921333, 24), to_signed(-1913928, 24), to_signed(-1906519, 24), to_signed(-1899105, 24), to_signed(-1891686, 24), to_signed(-1884263, 24), to_signed(-1876836, 24), to_signed(-1869404, 24), to_signed(-1861967, 24), to_signed(-1854527, 24), to_signed(-1847082, 24), to_signed(-1839633, 24), to_signed(-1832179, 24), to_signed(-1824721, 24), to_signed(-1817259, 24), to_signed(-1809792, 24), to_signed(-1802321, 24), to_signed(-1794846, 24), to_signed(-1787367, 24), to_signed(-1779883, 24), to_signed(-1772396, 24), to_signed(-1764904, 24), to_signed(-1757408, 24), to_signed(-1749908, 24), to_signed(-1742404, 24), to_signed(-1734895, 24), to_signed(-1727383, 24), to_signed(-1719866, 24), to_signed(-1712346, 24), to_signed(-1704821, 24), to_signed(-1697293, 24), to_signed(-1689760, 24), to_signed(-1682224, 24), to_signed(-1674683, 24), to_signed(-1667139, 24), to_signed(-1659590, 24), to_signed(-1652038, 24), to_signed(-1644482, 24), to_signed(-1636922, 24), to_signed(-1629358, 24), to_signed(-1621790, 24), to_signed(-1614219, 24), to_signed(-1606643, 24), to_signed(-1599064, 24), to_signed(-1591481, 24), to_signed(-1583895, 24), to_signed(-1576304, 24), to_signed(-1568710, 24), to_signed(-1561112, 24), to_signed(-1553511, 24), to_signed(-1545906, 24), to_signed(-1538297, 24), to_signed(-1530685, 24), to_signed(-1523069, 24), to_signed(-1515449, 24), to_signed(-1507826, 24), to_signed(-1500200, 24), to_signed(-1492570, 24), to_signed(-1484936, 24), to_signed(-1477299, 24), to_signed(-1469658, 24), to_signed(-1462014, 24), to_signed(-1454366, 24), to_signed(-1446715, 24), to_signed(-1439061, 24), to_signed(-1431403, 24), to_signed(-1423742, 24), to_signed(-1416078, 24), to_signed(-1408410, 24), to_signed(-1400739, 24), to_signed(-1393064, 24), to_signed(-1385387, 24), to_signed(-1377706, 24), to_signed(-1370021, 24), to_signed(-1362334, 24), to_signed(-1354643, 24), to_signed(-1346950, 24), to_signed(-1339253, 24), to_signed(-1331552, 24), to_signed(-1323849, 24), to_signed(-1316143, 24), to_signed(-1308433, 24), to_signed(-1300721, 24), to_signed(-1293005, 24), to_signed(-1285286, 24), to_signed(-1277565, 24), to_signed(-1269840, 24), to_signed(-1262112, 24), to_signed(-1254382, 24), to_signed(-1246648, 24), to_signed(-1238912, 24), to_signed(-1231172, 24), to_signed(-1223430, 24), to_signed(-1215685, 24), to_signed(-1207936, 24), to_signed(-1200186, 24), to_signed(-1192432, 24), to_signed(-1184675, 24), to_signed(-1176916, 24), to_signed(-1169154, 24), to_signed(-1161389, 24), to_signed(-1153621, 24), to_signed(-1145851, 24), to_signed(-1138078, 24), to_signed(-1130302, 24), to_signed(-1122524, 24), to_signed(-1114743, 24), to_signed(-1106959, 24), to_signed(-1099173, 24), to_signed(-1091384, 24), to_signed(-1083593, 24), to_signed(-1075799, 24), to_signed(-1068002, 24), to_signed(-1060204, 24), to_signed(-1052402, 24), to_signed(-1044598, 24), to_signed(-1036792, 24), to_signed(-1028983, 24), to_signed(-1021172, 24), to_signed(-1013358, 24), to_signed(-1005542, 24), to_signed(-997723, 24), to_signed(-989903, 24), to_signed(-982080, 24), to_signed(-974254, 24), to_signed(-966427, 24), to_signed(-958597, 24), to_signed(-950764, 24), to_signed(-942930, 24), to_signed(-935093, 24), to_signed(-927254, 24), to_signed(-919413, 24), to_signed(-911570, 24), to_signed(-903725, 24), to_signed(-895877, 24), to_signed(-888028, 24), to_signed(-880176, 24), to_signed(-872322, 24), to_signed(-864466, 24), to_signed(-856608, 24), to_signed(-848749, 24), to_signed(-840887, 24), to_signed(-833023, 24), to_signed(-825157, 24), to_signed(-817289, 24), to_signed(-809420, 24), to_signed(-801548, 24), to_signed(-793675, 24), to_signed(-785799, 24), to_signed(-777922, 24), to_signed(-770043, 24), to_signed(-762162, 24), to_signed(-754280, 24), to_signed(-746395, 24), to_signed(-738509, 24), to_signed(-730621, 24), to_signed(-722732, 24), to_signed(-714840, 24), to_signed(-706947, 24), to_signed(-699053, 24), to_signed(-691156, 24), to_signed(-683258, 24), to_signed(-675359, 24), to_signed(-667458, 24), to_signed(-659555, 24), to_signed(-651651, 24), to_signed(-643745, 24), to_signed(-635838, 24), to_signed(-627929, 24), to_signed(-620019, 24), to_signed(-612107, 24), to_signed(-604194, 24), to_signed(-596279, 24), to_signed(-588363, 24), to_signed(-580446, 24), to_signed(-572527, 24), to_signed(-564607, 24), to_signed(-556686, 24), to_signed(-548763, 24), to_signed(-540839, 24), to_signed(-532914, 24), to_signed(-524987, 24), to_signed(-517059, 24), to_signed(-509130, 24), to_signed(-501200, 24), to_signed(-493269, 24), to_signed(-485336, 24), to_signed(-477403, 24), to_signed(-469468, 24), to_signed(-461532, 24), to_signed(-453595, 24), to_signed(-445657, 24), to_signed(-437718, 24), to_signed(-429778, 24), to_signed(-421836, 24), to_signed(-413894, 24), to_signed(-405951, 24), to_signed(-398007, 24), to_signed(-390062, 24), to_signed(-382116, 24), to_signed(-374169, 24), to_signed(-366222, 24), to_signed(-358273, 24), to_signed(-350324, 24), to_signed(-342373, 24), to_signed(-334422, 24), to_signed(-326471, 24), to_signed(-318518, 24), to_signed(-310565, 24), to_signed(-302611, 24), to_signed(-294656, 24), to_signed(-286700, 24), to_signed(-278744, 24), to_signed(-270787, 24), to_signed(-262830, 24), to_signed(-254872, 24), to_signed(-246913, 24), to_signed(-238954, 24), to_signed(-230994, 24), to_signed(-223034, 24), to_signed(-215073, 24), to_signed(-207112, 24), to_signed(-199150, 24), to_signed(-191187, 24), to_signed(-183225, 24), to_signed(-175261, 24), to_signed(-167298, 24), to_signed(-159334, 24), to_signed(-151369, 24), to_signed(-143405, 24), to_signed(-135440, 24), to_signed(-127474, 24), to_signed(-119508, 24), to_signed(-111542, 24), to_signed(-103576, 24), to_signed(-95610, 24), to_signed(-87643, 24), to_signed(-79676, 24), to_signed(-71709, 24), to_signed(-63742, 24), to_signed(-55774, 24), to_signed(-47807, 24), to_signed(-39839, 24), to_signed(-31871, 24), to_signed(-23903, 24), to_signed(-15935, 24), to_signed(-7967, 24)
);
end sinewave;
