
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.fixed_pkg.ALL;
LIBRARY work;
USE work.arraypkg.all;
package mask_gen is
    CONSTANT decimal_numbers: mask := (
0 => to_sfixed(0.000000000000000000, mask_point'left, mask_point'right),
1 => to_sfixed(-0.000002997657576790, mask_point'left, mask_point'right),
2 => to_sfixed(-0.000032270637624758, mask_point'left, mask_point'right),
3 => to_sfixed(-0.000109196906789435, mask_point'left, mask_point'right),
4 => to_sfixed(-0.000229146304062663, mask_point'left, mask_point'right),
5 => to_sfixed(-0.000348429883709536, mask_point'left, mask_point'right),
6 => to_sfixed(-0.000382340622756462, mask_point'left, mask_point'right),
7 => to_sfixed(-0.000220615274892769, mask_point'left, mask_point'right),
8 => to_sfixed(0.000236695724375715, mask_point'left, mask_point'right),
9 => to_sfixed(0.001026777216200687, mask_point'left, mask_point'right),
10 => to_sfixed(0.002067851533207648, mask_point'left, mask_point'right),
11 => to_sfixed(0.003120191228069858, mask_point'left, mask_point'right),
12 => to_sfixed(0.003788488498053564, mask_point'left, mask_point'right),
13 => to_sfixed(0.003584529680295457, mask_point'left, mask_point'right),
14 => to_sfixed(0.002054436614102493, mask_point'left, mask_point'right),
15 => to_sfixed(-0.001046994209172248, mask_point'left, mask_point'right),
16 => to_sfixed(-0.005575114535046163, mask_point'left, mask_point'right),
17 => to_sfixed(-0.010863455454153802, mask_point'left, mask_point'right),
18 => to_sfixed(-0.015698258281229810, mask_point'left, mask_point'right),
19 => to_sfixed(-0.018439427364896319, mask_point'left, mask_point'right),
20 => to_sfixed(-0.017293417989963655, mask_point'left, mask_point'right),
21 => to_sfixed(-0.010699840337940400, mask_point'left, mask_point'right),
22 => to_sfixed(0.002247271459292921, mask_point'left, mask_point'right),
23 => to_sfixed(0.021447235827590182, mask_point'left, mask_point'right),
24 => to_sfixed(0.045611703314881916, mask_point'left, mask_point'right),
25 => to_sfixed(0.072326118112456927, mask_point'left, mask_point'right),
26 => to_sfixed(0.098370331720248047, mask_point'left, mask_point'right),
27 => to_sfixed(0.120250086520838281, mask_point'left, mask_point'right),
28 => to_sfixed(0.134833445023436971, mask_point'left, mask_point'right),
29 => to_sfixed(0.139952685973528335, mask_point'left, mask_point'right),
30 => to_sfixed(0.134833445023436999, mask_point'left, mask_point'right),
31 => to_sfixed(0.120250086520838281, mask_point'left, mask_point'right),
32 => to_sfixed(0.098370331720248047, mask_point'left, mask_point'right),
33 => to_sfixed(0.072326118112456914, mask_point'left, mask_point'right),
34 => to_sfixed(0.045611703314881909, mask_point'left, mask_point'right),
35 => to_sfixed(0.021447235827590193, mask_point'left, mask_point'right),
36 => to_sfixed(0.002247271459292922, mask_point'left, mask_point'right),
37 => to_sfixed(-0.010699840337940400, mask_point'left, mask_point'right),
38 => to_sfixed(-0.017293417989963658, mask_point'left, mask_point'right),
39 => to_sfixed(-0.018439427364896333, mask_point'left, mask_point'right),
40 => to_sfixed(-0.015698258281229820, mask_point'left, mask_point'right),
41 => to_sfixed(-0.010863455454153809, mask_point'left, mask_point'right),
42 => to_sfixed(-0.005575114535046163, mask_point'left, mask_point'right),
43 => to_sfixed(-0.001046994209172249, mask_point'left, mask_point'right),
44 => to_sfixed(0.002054436614102496, mask_point'left, mask_point'right),
45 => to_sfixed(0.003584529680295458, mask_point'left, mask_point'right),
46 => to_sfixed(0.003788488498053569, mask_point'left, mask_point'right),
47 => to_sfixed(0.003120191228069862, mask_point'left, mask_point'right),
48 => to_sfixed(0.002067851533207647, mask_point'left, mask_point'right),
49 => to_sfixed(0.001026777216200687, mask_point'left, mask_point'right),
50 => to_sfixed(0.000236695724375715, mask_point'left, mask_point'right),
51 => to_sfixed(-0.000220615274892769, mask_point'left, mask_point'right),
52 => to_sfixed(-0.000382340622756461, mask_point'left, mask_point'right),
53 => to_sfixed(-0.000348429883709536, mask_point'left, mask_point'right),
54 => to_sfixed(-0.000229146304062663, mask_point'left, mask_point'right),
55 => to_sfixed(-0.000109196906789435, mask_point'left, mask_point'right),
56 => to_sfixed(-0.000032270637624758, mask_point'left, mask_point'right),
57 => to_sfixed(-0.000002997657576790, mask_point'left, mask_point'right),
58 => to_sfixed(0.000000000000000000, mask_point'left, mask_point'right)

);
END mask_gen;
